module prefix_decode (
       	mask_prefix,
        pre_seg_override,
        pre_seg_override_valid,
        pre_repeat,
        pre_size_override			
);

  input [23:0]      mask_prefix;
  output [2:0]      pre_seg_override;
  output            pre_seg_override_valid;
  output            pre_repeat;
  output            pre_size_override;


   assign i23 = mask_prefix[23];
   assign i22 = mask_prefix[22];
   assign i21 = mask_prefix[21];
   assign i20 = mask_prefix[20];
   assign i19 = mask_prefix[19];
   assign i18 = mask_prefix[18];
   assign i17 = mask_prefix[17];
   assign i16 = mask_prefix[16];
   assign i15 = mask_prefix[15];
   assign i14 = mask_prefix[14];
   assign i13 = mask_prefix[13];
   assign i12 = mask_prefix[12];
   assign i11 = mask_prefix[11];
   assign i10 = mask_prefix[10];
   assign i9 = mask_prefix[9];
   assign i8 = mask_prefix[8];
   assign i7 = mask_prefix[7];
   assign i6 = mask_prefix[6];
   assign i5 = mask_prefix[5];
   assign i4 = mask_prefix[4];
   assign i3 = mask_prefix[3];
   assign i2 = mask_prefix[2];
   assign i1 = mask_prefix[1];
   assign i0 = mask_prefix[0];  
   
wire i23_not;
wire i22_not;
wire i19_not;
wire i18_not;
wire i17_not;
wire i16_not;
wire i15_not;
wire i14_not;
wire i13_not;
wire i11_not;
wire i10_not;
wire i7_not;
wire i2_not;
wire i1_not;
wire and0;
wire i22_not;
wire i14_not;
wire and1;
wire i21_not;
wire i20_not;
wire i12_not;
wire i9_not;
wire i6_not;
wire i5_not;
wire and2;
wire i5_not;
wire and3;
wire i13_not;
wire i8_not;
wire i4_not;
wire i0_not;
wire and4;
wire i3_not;
wire and5;
wire and6;
wire i3_not;
wire i2_not;
wire and7;
wire and8;
wire i18_not;
wire i1_not;
wire and9;
wire and10;
wire and11;
wire i23_not;
wire i8_not;
wire and12;
wire and13;
wire and14;
wire and15;
wire and16;
wire and17;
wire and18;
wire and19;
wire and20;
wire and21;
wire and22;
wire and23;
wire and24;
wire i20_not;
wire and25;
wire i7_not;
wire and26;
wire and27;
wire and28;
wire i11_not;
wire and29;
wire and30;
wire and31;
wire and32;
wire i20_not;
wire and33;
wire and34;
wire and35;
wire and36;
wire and37;
wire or0;
wire i12_not;
wire and38;
wire and39;
wire and40;
wire and41;
wire and42;
wire and43;
wire and44;
wire i16_not;
wire and45;
wire and46;
wire and47;
wire and48;
wire and49;
wire i21_not;
wire and50;
wire and51;
wire i19_not;
wire and52;
wire and53;
wire and54;
wire and55;
wire and56;
wire and57;
wire and58;
wire and59;
wire and60;
wire i6_not;
wire and61;
wire and62;
wire i10_not;
wire and63;
wire and64;
wire and65;
wire and66;
wire and67;
wire and68;
wire and69;
wire and70;
wire and71;
wire and72;
wire and73;
wire and74;
wire i8_not;
wire and75;
wire and76;
wire or1;
wire and77;
wire and78;
wire and79;
wire and80;
wire and81;
wire and82;
wire and83;
wire and84;
wire and85;
wire and86;
wire and87;
wire and88;
wire and89;
wire and90;
wire and91;
wire and92;
wire and93;
wire and94;
wire and95;
wire and96;
wire and97;
wire i17_not;
wire and98;
wire and99;
wire and100;
wire and101;
wire and102;
wire and103;
wire and104;
wire and105;
wire and106;
wire and107;
wire and108;
wire and109;
wire or2;
wire and110;
wire and111;
wire and112;
wire and113;
wire and114;
wire i15_not;
wire and115;
wire and116;
wire and117;
wire and118;
wire and119;
wire and120;
wire and121;
wire and122;
wire and123;
wire and124;
wire and125;
wire and126;
wire i4_not;
wire and127;
wire and128;
wire and129;
wire and130;
wire and131;
wire and132;
wire and133;
wire and134;
wire and135;
wire and136;
wire and137;
wire i11_not;
wire and138;
wire and139;
wire and140;
wire and141;
wire or3;
wire and142;
wire i17_not;
wire and143;
wire and144;
wire and145;
wire and146;
wire and147;
wire i23_not;
wire and148;
wire and149;
wire and150;
wire and151;
wire and152;
wire and153;
wire and154;
wire and155;
wire and156;
wire and157;
wire and158;
wire and159;
wire and160;
wire and161;
wire and162;
wire and163;
wire and164;
wire and165;
wire and166;
wire and167;
wire and168;
wire and169;
wire and170;
wire and171;
wire and172;
wire and173;
wire or4;
wire and174;
wire and175;
wire and176;
wire and177;
wire and178;
wire and179;
wire and180;
wire and181;
wire and182;
wire and183;
wire and184;
wire and185;
wire and186;
wire and187;
wire and188;
wire and189;
wire and190;
wire and191;
wire and192;
wire and193;
wire and194;
wire and195;
wire and196;
wire and197;
wire and198;
wire and199;
wire and200;
wire and201;
wire and202;
wire and203;
wire or5;

inv1$ i22_inv (.out(i22_not), .in(i22));
inv1$ i19_inv (.out(i19_not), .in(i19));
inv1$ i18_inv (.out(i18_not), .in(i18));
inv1$ i17_inv (.out(i17_not), .in(i17));
inv1$ i16_inv (.out(i16_not), .in(i16));
inv1$ i15_inv (.out(i15_not), .in(i15));
inv1$ i14_inv (.out(i14_not), .in(i14));
inv1$ i13_inv (.out(i13_not), .in(i13));
inv1$ i11_inv (.out(i11_not), .in(i11));
inv1$ i10_inv (.out(i10_not), .in(i10));
inv1$ i7_inv (.out(i7_not), .in(i7));
inv1$ i2_inv (.out(i2_not), .in(i2));
inv1$ i1_inv (.out(i1_not), .in(i1));
inv1$ i21_inv (.out(i21_not), .in(i21));
inv1$ i20_inv (.out(i20_not), .in(i20));
inv1$ i12_inv (.out(i12_not), .in(i12));
inv1$ i9_inv (.out(i9_not), .in(i9));
inv1$ i6_inv (.out(i6_not), .in(i6));
inv1$ i5_inv (.out(i5_not), .in(i5));
inv1$ i8_inv (.out(i8_not), .in(i8));
inv1$ i4_inv (.out(i4_not), .in(i4));
inv1$ i0_inv (.out(i0_not), .in(i0));
inv1$ i23_inv (.out(i23_not), .in(i23));

and24$ and_gate0(.out(and0), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17_not), .in7(i16_not), .in8(i15_not), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11_not), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate1(.out(and1), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15_not), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6
), .in18(i5), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate2(.out(and2), .in0(i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17), .in7(i16), .in8(i15), .in9(i14
), .in10(i13_not), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate3(.out(and3), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16_not), .in8(i15), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate4(.out(and4), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate5(.out(and5), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20
), .in4(i19), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0_not));
and24$ and_gate6(.out(and6), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16_not), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12
), .in12(i11_not), .in13(i10_not), .in14(i9), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate7(.out(and7), .in0(i23), .in1(i22_not), .in2(i21_not), .in3(i20), .in4(i19
), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7_not), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate8(.out(and8), .in0(i23), .in1(i22_not), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11
), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate9(.out(and9), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate10(.out(and10), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14), .in10(i13_not), .in11(i12_not), .in12(i11), .in13(i10
), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate11(.out(and11), .in0(i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17
), .in7(i16_not), .in8(i15), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate12(.out(and12), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate13(.out(and13), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16
), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0));
and24$ and_gate14(.out(and14), .in0(
i23), .in1(i22_not), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10_not), .in14(i9), .in15(i8
), .in16(i7_not), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate15(.out(and15), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18), .in6(i17), .in7(i16
), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate16(.out(and16), .in0(
i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7
), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0));
and24$ and_gate17(.out(and17), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16), .in8(i15
), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate18(.out(and18), .in0(i23), .in1(i22_not), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9), .in15(i8), .in16(i7), .in17(i6), .in18(i5
), .in19(i4_not), .in20(i3_not), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate19(.out(and19), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14
), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4), .in20(i3), .in21(i2), .in22(i1), .in23(i0));
and24$ and_gate20(.out(and20), .in0(i23_not), .in1(i22), .in2(i21
), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5), .in19(i4
), .in20(i3), .in21(i2), .in22(i1), .in23(i0));
and24$ and_gate21(.out(and21), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16_not), .in8(i15), .in9(i14), .in10(i13), .in11(i12
), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0_not));
and24$ and_gate22(.out(and22), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20
), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7), .in17(i6), .in18(i5), .in19(i4), .in20(i3), .in21(i2
), .in22(i1_not), .in23(i0_not));
and24$ and_gate23(.out(and23), .in0(i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11
), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate24(.out(and24), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18
), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and21$ and_gate25(.out(and25), .in0(i20_not), .in1(i19), .in2(i18_not), .in3(i17), .in4(i16_not), .in5(i15), .in6(i14), .in7(i13_not), .in8(i12), .in9(i11), .in10(i10), .in11(i9), .in12(i8), .in13(i7_not), .in14(i6_not), .in15(i5), .in16(i4
), .in17(i3_not), .in18(i2_not), .in19(i1), .in20(i0));
and18$ and_gate26(.out(and26), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13_not), .in5(i12_not), .in6(i11_not), .in7(i10_not), .in8(i9), .in9(i8_not), .in10(i7_not), .in11(i6), .in12(i5_not), .in13(i4_not), .in14(i3), .in15(i2), .in16(i1_not), .in17(i0));
and18$ and_gate27(.out(and27), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13_not), .in5(i12), .in6(i11_not), .in7(i10_not), .in8(i9
), .in9(i8_not), .in10(i7_not), .in11(i6), .in12(i5), .in13(i4_not), .in14(i3), .in15(i2), .in16(i1_not), .in17(i0));
and18$ and_gate28(.out(and28), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13), .in5(i12_not), .in6(i11
), .in7(i10_not), .in8(i9), .in9(i8_not), .in10(i7), .in11(i6), .in12(i5_not), .in13(i4_not), .in14(i3), .in15(i2_not), .in16(i1), .in17(i0));
and16$ and_gate29(.out(and29), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i11_not), .in5(i10), .in6(i9_not), .in7(i8), .in8(i7_not), .in9(i6_not), .in10(i5_not), .in11(i4_not), .in12(i3), .in13(i2), .in14(i1), .in15(i0));
and16$ and_gate30(.out(and30), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19), .in5(i18
), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14), .in10(i5_not), .in11(i4), .in12(i3_not), .in13(i2), .in14(i1_not), .in15(i0));
and16$ and_gate31(.out(and31), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18
), .in6(i17_not), .in7(i8_not), .in8(i7), .in9(i6_not), .in10(i5), .in11(i4_not), .in12(i3_not), .in13(i2), .in14(i1_not), .in15(i0));
and16$ and_gate32(.out(and32), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and16$ and_gate33(.out(and33), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i8_not), .in8(i7), .in9(i6_not), .in10(i5), .in11(i4_not), .in12(i3_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and16$ and_gate34(.out(and34), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and16$ and_gate35(.out(and35), .in0(i23), .in1(i22), .in2(i21
), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and16$ and_gate36(.out(and36), .in0(i23), .in1(i22
), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14_not), .in10(i5_not), .in11(i4), .in12(i3_not), .in13(i2), .in14(i1_not), .in15(i0_not));
and9$ and_gate37(.out(and37), .in0(i8_not), .in1(i7_not), .in2(i6), .in3(i5_not), .in4(i4_not), .in5(i3_not), .in6(i2_not), .in7(i1), .in8(i0_not));
and24$ and_gate38(.out(and38), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14), .in10(i13_not), .in11(i12_not), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate39(.out(and39), .in0(i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate40(.out(and40), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate41(.out(and41), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18
), .in6(i17), .in7(i16_not), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate42(.out(and42), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10
), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate43(.out(and43), .in0(i23), .in1(i22), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17
), .in7(i16), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7_not), .in17(i6_not), .in18(i5), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate44(.out(and44), .in0(
i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8
), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate45(.out(and45), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate46(.out(and46), .in0(
i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7
), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0));
and24$ and_gate47(.out(and47), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16), .in8(i15
), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate48(.out(and48), .in0(i23), .in1(i22_not), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9), .in15(i8), .in16(i7), .in17(i6), .in18(i5
), .in19(i4_not), .in20(i3_not), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate49(.out(and49), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14
), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3_not), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate50(.out(and50), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16_not), .in8(i15), .in9(i14), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5), .in19(i4
), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0_not));
and23$ and_gate51(.out(and51), .in0(i23), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18), .in6(i16), .in7(i15), .in8(i14), .in9(i13_not), .in10(i12_not), .in11(i11), .in12(i10), .in13(i9_not), .in14(i8_not), .in15(i7), .in16(i6), .in17(i5_not), .in18(i4), .in19(i3), .in20(i2), .in21(i1), .in22(i0_not));
and24$ and_gate52(.out(and52), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7), .in17(i6), .in18(i5), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate53(.out(and53), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1), .in23(i0_not));
and23$ and_gate54(.out(and54), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i19), .in4(i18), .in5(i17
), .in6(i16_not), .in7(i15), .in8(i14), .in9(i13), .in10(i12), .in11(i11_not), .in12(i10_not), .in13(i9), .in14(i8), .in15(i7_not), .in16(i6), .in17(i5), .in18(i4_not), .in19(i3_not), .in20(i2), .in21(i1), .in22(i0_not));
and24$ and_gate55(.out(and55), .in0(
i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and21$ and_gate56(.out(and56), .in0(i20_not), .in1(i19), .in2(i18_not), .in3(i17), .in4(i16_not), .in5(i15), .in6(i14_not), .in7(i13
), .in8(i12_not), .in9(i11_not), .in10(i10_not), .in11(i9), .in12(i8), .in13(i7_not), .in14(i6), .in15(i5), .in16(i4_not), .in17(i3_not), .in18(i2), .in19(i1), .in20(i0_not));
and21$ and_gate57(.out(and57), .in0(i20_not), .in1(i19), .in2(i18_not), .in3(i17), .in4(i16_not), .in5(i15_not), .in6(i14_not), .in7(i13), .in8(i12_not), .in9(i11_not), .in10(i10_not), .in11(i9), .in12(i8_not), .in13(i7_not), .in14(i6), .in15(i5), .in16(i4_not), .in17(i3_not), .in18(i2), .in19(i1
), .in20(i0_not));
and24$ and_gate58(.out(and58), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10
), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and21$ and_gate59(.out(and59), .in0(i20_not), .in1(i19), .in2(i18_not), .in3(i17), .in4(i16), .in5(i15_not), .in6(i14
), .in7(i13), .in8(i12_not), .in9(i11_not), .in10(i10), .in11(i9), .in12(i8_not), .in13(i7_not), .in14(i6), .in15(i5_not), .in16(i4), .in17(i3_not), .in18(i2), .in19(i1), .in20(i0_not));
and21$ and_gate60(.out(and60), .in0(i20_not), .in1(i19
), .in2(i18_not), .in3(i17), .in4(i16), .in5(i15_not), .in6(i14), .in7(i13), .in8(i12_not), .in9(i11), .in10(i10), .in11(i9), .in12(i8), .in13(i7_not), .in14(i6_not), .in15(i5), .in16(i4), .in17(i3_not), .in18(i2), .in19(i1
), .in20(i0_not));
and21$ and_gate61(.out(and61), .in0(i20_not), .in1(i19), .in2(i18_not), .in3(i17), .in4(i16_not), .in5(i15), .in6(i14), .in7(i13_not), .in8(i12), .in9(i11), .in10(i10), .in11(i9), .in12(i8), .in13(i7_not), .in14(i6_not), .in15(i5), .in16(i4), .in17(i3_not), .in18(i2_not), .in19(i1), .in20(i0));
and18$ and_gate62(.out(and62), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13_not), .in5(i12_not), .in6(i11_not), .in7(i10_not), .in8(i9), .in9(i8_not), .in10(i7_not), .in11(i6), .in12(i5_not), .in13(i4_not), .in14(i3), .in15(i2), .in16(i1_not), .in17(i0));
and18$ and_gate63(.out(and63), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13_not), .in5(i12), .in6(i11_not), .in7(i10_not), .in8(i9), .in9(i8_not), .in10(i7_not), .in11(i6), .in12(i5), .in13(i4_not), .in14(i3), .in15(i2), .in16(i1_not), .in17(i0));
and18$ and_gate64(.out(and64), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13), .in5(i12_not), .in6(i11
), .in7(i10_not), .in8(i9), .in9(i8_not), .in10(i7), .in11(i6), .in12(i5_not), .in13(i4_not), .in14(i3), .in15(i2_not), .in16(i1), .in17(i0));
and18$ and_gate65(.out(and65), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13_not), .in5(i12), .in6(i11), .in7(i10), .in8(i9_not), .in9(i8), .in10(i7), .in11(i6), .in12(i5), .in13(i4_not), .in14(i3_not), .in15(i2), .in16(i1), .in17(i0_not));
and16$ and_gate66(.out(and66), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20
), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14), .in10(i5_not), .in11(i4), .in12(i3_not), .in13(i2), .in14(i1_not), .in15(i0));
and16$ and_gate67(.out(and67), .in0(i23), .in1(i22), .in2(i21), .in3(i20
), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9_not), .in15(i8_not));
and16$ and_gate68(.out(and68), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14), .in10(i5_not), .in11(i4), .in12(i3_not), .in13(i2), .in14(i1), .in15(i0_not));
and16$ and_gate69(.out(and69), .in0(i23_not), .in1(i22
), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18), .in6(i17_not), .in7(i8_not), .in8(i7), .in9(i6_not), .in10(i5), .in11(i4_not), .in12(i3_not), .in13(i2), .in14(i1_not), .in15(i0));
and16$ and_gate70(.out(and70), .in0(i23_not), .in1(i22
), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not));
and16$ and_gate71(.out(and71), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and16$ and_gate72(.out(and72), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i8_not), .in8(i7), .in9(i6_not), .in10(i5), .in11(i4_not), .in12(i3_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and16$ and_gate73(.out(and73), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and16$ and_gate74(.out(and74), .in0(
i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14_not), .in10(i5_not), .in11(i4), .in12(i3_not), .in13(i2), .in14(i1_not), .in15(i0_not));
and9$ and_gate75(.out(and75), .in0(i8_not), .in1(i7_not), .in2(i6), .in3(i5), .in4(i4), .in5(i3_not), .in6(i2_not), .in7(i1_not), .in8(i0_not));
and9$ and_gate76(.out(and76), .in0(i8_not), .in1(i7_not), .in2(i6), .in3(i5_not), .in4(i4_not), .in5(i3_not), .in6(i2_not), .in7(i1), .in8(i0_not));
and24$ and_gate77(.out(and77), .in0(i23), .in1(i22), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate78(.out(and78), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19
), .in5(i18), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6_not), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate79(.out(and79), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14), .in10(i13_not), .in11(i12_not), .in12(i11
), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate80(.out(and80), .in0(i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19
), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1
), .in23(i0));
and24$ and_gate81(.out(and81), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10
), .in14(i9), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate82(.out(and82), .in0(i23), .in1(i22), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17
), .in7(i16), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7_not), .in17(i6_not), .in18(i5), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate83(.out(and83), .in0(
i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8
), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate84(.out(and84), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate85(.out(and85), .in0(
i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7
), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0));
and24$ and_gate86(.out(and86), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15
), .in9(i14), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3_not), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate87(.out(and87), .in0(i23_not), .in1(i22
), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16_not), .in8(i15), .in9(i14), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5
), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0_not));
and23$ and_gate88(.out(and88), .in0(i23), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18), .in6(i16), .in7(i15), .in8(i14), .in9(i13_not), .in10(i12_not), .in11(i11), .in12(i10), .in13(i9_not), .in14(i8_not), .in15(i7), .in16(i6), .in17(i5_not), .in18(i4), .in19(i3), .in20(i2), .in21(i1), .in22(i0_not));
and24$ and_gate89(.out(and89), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19
), .in5(i18), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1
), .in23(i0));
and24$ and_gate90(.out(and90), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10
), .in14(i9), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1), .in23(i0_not));
and23$ and_gate91(.out(and91), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i19), .in4(i18), .in5(i17), .in6(i16_not), .in7(i15), .in8(i14), .in9(i13), .in10(i12), .in11(i11_not), .in12(i10_not), .in13(i9), .in14(i8), .in15(i7_not), .in16(i6), .in17(i5), .in18(i4_not), .in19(i3_not), .in20(i2), .in21(i1), .in22(i0_not));
and24$ and_gate92(.out(and92), .in0(i23
), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7
), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and21$ and_gate93(.out(and93), .in0(i20_not), .in1(i19), .in2(i18_not), .in3(i17), .in4(i16_not), .in5(i15), .in6(i14_not), .in7(i13), .in8(i12_not), .in9(i11_not), .in10(i10_not), .in11(i9), .in12(i8), .in13(i7_not), .in14(i6), .in15(i5), .in16(i4_not), .in17(i3_not), .in18(i2), .in19(i1), .in20(i0_not));
and21$ and_gate94(.out(and94), .in0(i20_not), .in1(i19), .in2(i18_not), .in3(i17
), .in4(i16_not), .in5(i15_not), .in6(i14_not), .in7(i13), .in8(i12_not), .in9(i11_not), .in10(i10_not), .in11(i9), .in12(i8_not), .in13(i7_not), .in14(i6), .in15(i5), .in16(i4_not), .in17(i3_not), .in18(i2), .in19(i1), .in20(i0_not));
and24$ and_gate95(.out(and95), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and21$ and_gate96(.out(and96), .in0(i20_not), .in1(i19), .in2(i18_not), .in3(i17), .in4(i16), .in5(i15_not), .in6(i14), .in7(i13), .in8(i12_not), .in9(i11_not), .in10(i10), .in11(i9), .in12(i8_not), .in13(i7_not), .in14(i6), .in15(i5_not), .in16(i4), .in17(i3_not), .in18(i2), .in19(i1), .in20(i0_not));
and21$ and_gate97(.out(and97), .in0(i20_not), .in1(i19), .in2(i18_not), .in3(i17
), .in4(i16_not), .in5(i15), .in6(i14), .in7(i13_not), .in8(i12), .in9(i11), .in10(i10), .in11(i9), .in12(i8), .in13(i7_not), .in14(i6_not), .in15(i5), .in16(i4), .in17(i3_not), .in18(i2_not), .in19(i1), .in20(i0));
and18$ and_gate98(.out(and98), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13_not), .in5(i12_not), .in6(i11_not), .in7(i10_not), .in8(i9), .in9(i8_not), .in10(i7_not), .in11(i6), .in12(i5_not), .in13(i4_not), .in14(i3), .in15(i2), .in16(i1_not), .in17(i0));
and18$ and_gate99(.out(and99), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13_not), .in5(i12), .in6(i11_not), .in7(i10_not), .in8(i9), .in9(i8_not), .in10(i7_not), .in11(i6), .in12(i5), .in13(i4_not), .in14(i3
), .in15(i2), .in16(i1_not), .in17(i0));
and18$ and_gate100(.out(and100), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13), .in5(i12_not), .in6(i11), .in7(i10_not), .in8(i9), .in9(i8_not), .in10(i7), .in11(i6), .in12(i5_not), .in13(i4_not), .in14(i3), .in15(i2_not), .in16(i1), .in17(i0));
and18$ and_gate101(.out(and101), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13_not), .in5(i12), .in6(i11), .in7(i10), .in8(i9_not), .in9(i8), .in10(i7), .in11(i6
), .in12(i5), .in13(i4_not), .in14(i3_not), .in15(i2), .in16(i1), .in17(i0_not));
and16$ and_gate102(.out(and102), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18), .in6(i17_not), .in7(i8_not), .in8(i7), .in9(i6_not), .in10(i5), .in11(i4_not), .in12(i3_not), .in13(i2), .in14(i1_not), .in15(i0));
and16$ and_gate103(.out(and103), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i8_not), .in8(i7), .in9(i6_not), .in10(i5), .in11(i4_not), .in12(i3_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and16$ and_gate104(.out(and104), .in0(i23), .in1(i22), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and12$ and_gate105(.out(and105), .in0(i11_not), .in1(i10_not), .in2(i9), .in3(i8_not), .in4(i7_not), .in5(i6_not), .in6(i5_not), .in7(i4_not), .in8(i3), .in9(i2_not), .in10(i1), .in11(i0));
and9$ and_gate106(.out(and106), .in0(i8_not), .in1(i7_not), .in2(i6), .in3(i5), .in4(i4), .in5(i3_not), .in6(i2_not), .in7(i1_not), .in8(i0_not));
and8$ and_gate107(.out(and107), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17), .in7(i16_not));
and9$ and_gate108(.out(and108), .in0(i8_not), .in1(i7_not), .in2(i6), .in3(i5), .in4(i4_not), .in5(i3), .in6(i2), .in7(i1_not), .in8(i0_not));
and9$ and_gate109(.out(and109), .in0(i8_not), .in1(i7_not), .in2(i6
), .in3(i5_not), .in4(i4_not), .in5(i3_not), .in6(i2_not), .in7(i1), .in8(i0_not));
and24$ and_gate110(.out(and110), .in0(i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17), .in7(i16), .in8(i15), .in9(i14), .in10(i13_not), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate111(.out(and111), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1
), .in23(i0));
and24$ and_gate112(.out(and112), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate113(.out(and113), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14), .in10(i13_not), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate114(.out(and114), .in0(
i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8
), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate115(.out(and115), .in0(i23), .in1(i22), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7_not), .in17(i6_not), .in18(i5), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate116(.out(and116), .in0(i23), .in1(i22
), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate117(.out(and117), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0));
and24$ and_gate118(.out(and118), .in0(i23), .in1(i22_not), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6_not), .in18(i5), .in19(i4
), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate119(.out(and119), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18), .in6(i17), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate120(.out(and120), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3
), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate121(.out(and121), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14), .in10(i13), .in11(i12
), .in12(i11_not), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3_not), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate122(.out(and122), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4), .in20(i3), .in21(i2
), .in22(i1), .in23(i0));
and24$ and_gate123(.out(and123), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3), .in21(i2), .in22(i1), .in23(i0));
and24$ and_gate124(.out(and124), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16_not), .in8(i15), .in9(i14), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0_not));
and24$ and_gate125(.out(and125), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1), .in23(i0));
and24$ and_gate126(.out(and126), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7), .in17(i6), .in18(i5), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and23$ and_gate127(.out(and127), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i19), .in4(i18), .in5(i17), .in6(i16_not), .in7(i15), .in8(i14), .in9(i13), .in10(i12), .in11(i11_not), .in12(i10_not), .in13(i9), .in14(i8), .in15(i7_not), .in16(i6), .in17(i5), .in18(i4_not), .in19(i3_not), .in20(i2), .in21(i1), .in22(i0_not));
and24$ and_gate128(.out(and128), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13
), .in11(i12), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and21$ and_gate129(.out(and129), .in0(i20_not), .in1(i19), .in2(i18_not), .in3(i17
), .in4(i16), .in5(i15_not), .in6(i14), .in7(i13), .in8(i12_not), .in9(i11), .in10(i10), .in11(i9), .in12(i8), .in13(i7_not), .in14(i6_not), .in15(i5), .in16(i4), .in17(i3_not), .in18(i2), .in19(i1), .in20(i0_not));
and16$ and_gate130(.out(and130), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i11_not), .in5(i10), .in6(i9_not), .in7(i8), .in8(i7_not), .in9(i6_not), .in10(i5_not), .in11(i4_not), .in12(i3), .in13(i2), .in14(i1), .in15(i0));
and18$ and_gate131(.out(and131), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13_not), .in5(i12), .in6(i11), .in7(i10), .in8(i9_not), .in9(i8), .in10(i7), .in11(i6), .in12(i5), .in13(i4_not), .in14(i3_not), .in15(i2), .in16(i1), .in17(i0_not));
and16$ and_gate132(.out(and132), .in0(
i23), .in1(i22), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9_not), .in15(i8_not));
and16$ and_gate133(.out(and133), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18), .in6(i17_not), .in7(i8_not), .in8(i7), .in9(i6_not), .in10(i5), .in11(i4_not), .in12(i3_not), .in13(i2), .in14(i1_not), .in15(i0));
and16$ and_gate134(.out(and134), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not));
and16$ and_gate135(.out(and135), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i8_not), .in8(i7), .in9(i6_not), .in10(i5), .in11(i4_not), .in12(i3_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and16$ and_gate136(.out(and136), .in0(
i23), .in1(i22), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and16$ and_gate137(.out(and137), .in0(
i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14_not), .in10(i5_not), .in11(i4), .in12(i3_not), .in13(i2), .in14(i1_not), .in15(i0_not));
and12$ and_gate138(.out(and138), .in0(i11_not), .in1(i10_not), .in2(i9), .in3(i8_not), .in4(i7_not), .in5(i6_not), .in6(i5_not), .in7(i4_not), .in8(i3), .in9(i2_not), .in10(i1), .in11(i0));
and8$ and_gate139(.out(and139), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17), .in7(i16_not));
and9$ and_gate140(.out(and140), .in0(i8_not), .in1(i7_not), .in2(i6), .in3(i5), .in4(i4_not), .in5(i3), .in6(i2), .in7(i1_not), .in8(i0_not));
and9$ and_gate141(.out(and141), .in0(i8_not), .in1(i7_not), .in2(i6
), .in3(i5_not), .in4(i4_not), .in5(i3_not), .in6(i2_not), .in7(i1), .in8(i0_not));
and24$ and_gate142(.out(and142), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate143(.out(and143), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14), .in10(i13_not), .in11(i12_not), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate144(.out(and144), .in0(
i23), .in1(i22_not), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10_not), .in14(i9_not), .in15(i8
), .in16(i7_not), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate145(.out(and145), .in0(i23), .in1(i22_not), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18), .in6(i17), .in7(i16
), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate146(.out(and146), .in0(i23
), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8_not), .in16(i7
), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate147(.out(and147), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15
), .in9(i14), .in10(i13_not), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate148(.out(and148), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7
), .in17(i6_not), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate149(.out(and149), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2_not), .in22(i1_not), .in23(i0));
and24$ and_gate150(.out(and150), .in0(i23), .in1(i22
), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate151(.out(and151), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0));
and24$ and_gate152(.out(and152), .in0(i23_not), .in1(i22), .in2(i21
), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate153(.out(and153), .in0(i23), .in1(i22_not), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15_not), .in9(i14), .in10(i13
), .in11(i12), .in12(i11_not), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate154(.out(and154), .in0(i23_not), .in1(i22_not), .in2(i21
), .in3(i20), .in4(i19_not), .in5(i18), .in6(i17), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4
), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate155(.out(and155), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate156(.out(and156), .in0(i23), .in1(i22_not), .in2(i21_not), .in3(i20
), .in4(i19), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9), .in15(i8), .in16(i7), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3_not), .in21(i2
), .in22(i1), .in23(i0_not));
and24$ and_gate157(.out(and157), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3_not), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate158(.out(and158), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4), .in20(i3), .in21(i2), .in22(i1
), .in23(i0));
and24$ and_gate159(.out(and159), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10
), .in14(i9), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3), .in21(i2), .in22(i1), .in23(i0));
and24$ and_gate160(.out(and160), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17
), .in7(i16_not), .in8(i15), .in9(i14), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0_not));
and23$ and_gate161(.out(and161), .in0(
i23), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18), .in6(i16), .in7(i15), .in8(i14), .in9(i13_not), .in10(i12_not), .in11(i11), .in12(i10), .in13(i9_not), .in14(i8_not), .in15(i7), .in16(i6
), .in17(i5_not), .in18(i4), .in19(i3), .in20(i2), .in21(i1), .in22(i0_not));
and24$ and_gate162(.out(and162), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7), .in17(i6), .in18(i5), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate163(.out(and163), .in0(i23_not), .in1(i22_not), .in2(i21
), .in3(i20), .in4(i19), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4
), .in20(i3), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate164(.out(and164), .in0(i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13), .in11(i12
), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and19$ and_gate165(.out(and165), .in0(i23), .in1(i22_not), .in2(i21_not), .in3(i20_not), .in4(i19_not), .in5(i18), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7_not), .in17(i6), .in18(i5));
and19$ and_gate166(.out(and166), .in0(i23
), .in1(i22), .in2(i21), .in3(i20), .in4(i19), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7), .in17(i6
), .in18(i5_not));
and21$ and_gate167(.out(and167), .in0(i20_not), .in1(i19), .in2(i18_not), .in3(i17), .in4(i16_not), .in5(i15), .in6(i14), .in7(i13_not), .in8(i12), .in9(i11), .in10(i10), .in11(i9), .in12(i8), .in13(i7_not), .in14(i6_not), .in15(i5), .in16(i4), .in17(i3_not), .in18(i2_not), .in19(i1), .in20(i0));
and16$ and_gate168(.out(and168), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i11_not), .in5(i10), .in6(i9_not), .in7(i8), .in8(i7_not), .in9(i6_not), .in10(i5_not), .in11(i4_not), .in12(i3), .in13(i2), .in14(i1), .in15(i0));
and18$ and_gate169(.out(and169), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13_not), .in5(i12), .in6(i11), .in7(i10), .in8(i9_not), .in9(i8), .in10(i7), .in11(i6
), .in12(i5), .in13(i4_not), .in14(i3_not), .in15(i2), .in16(i1), .in17(i0_not));
and16$ and_gate170(.out(and170), .in0(i23), .in1(i22), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14
), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9_not), .in15(i8_not));
and16$ and_gate171(.out(and171), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14), .in10(i5_not), .in11(i4), .in12(i3_not), .in13(i2), .in14(i1), .in15(i0_not));
and16$ and_gate172(.out(and172), .in0(i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16
), .in8(i15), .in9(i14_not), .in10(i5_not), .in11(i4), .in12(i3_not), .in13(i2), .in14(i1_not), .in15(i0_not));
and9$ and_gate173(.out(and173), .in0(i8_not), .in1(i7_not), .in2(i6), .in3(i5), .in4(i4_not), .in5(i3), .in6(i2), .in7(i1_not), .in8(i0_not));
and24$ and_gate174(.out(and174), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15), .in9(i14), .in10(i13), .in11(i12
), .in12(i11_not), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3_not), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate175(.out(and175), .in0(i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19
), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14), .in10(i13_not), .in11(i12_not), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2
), .in22(i1_not), .in23(i0_not));
and24$ and_gate176(.out(and176), .in0(i23), .in1(i22_not), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7_not), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate177(.out(and177), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19
), .in5(i18), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate178(.out(and178), .in0(i23_not), .in1(i22), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11
), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and24$ and_gate179(.out(and179), .in0(i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19
), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7), .in17(i6_not), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2
), .in22(i1_not), .in23(i0_not));
and24$ and_gate180(.out(and180), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate181(.out(and181), .in0(i23), .in1(i22_not), .in2(i21_not), .in3(i20), .in4(i19
), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10_not), .in14(i9), .in15(i8), .in16(i7_not), .in17(i6_not), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate182(.out(and182), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18), .in6(i17), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13_not), .in11(i12), .in12(i11
), .in13(i10_not), .in14(i9_not), .in15(i8), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4), .in20(i3_not), .in21(i2_not), .in22(i1), .in23(i0));
and24$ and_gate183(.out(and183), .in0(i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18
), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13_not), .in11(i12), .in12(i11), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0));
and24$ and_gate184(.out(and184), .in0(
i23), .in1(i22_not), .in2(i21_not), .in3(i20), .in4(i19), .in5(i18_not), .in6(i17_not), .in7(i16), .in8(i15), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11), .in13(i10), .in14(i9), .in15(i8), .in16(i7
), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3_not), .in21(i2), .in22(i1), .in23(i0_not));
and23$ and_gate185(.out(and185), .in0(i23), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18), .in6(i16), .in7(i15), .in8(i14
), .in9(i13_not), .in10(i12_not), .in11(i11), .in12(i10), .in13(i9_not), .in14(i8_not), .in15(i7), .in16(i6), .in17(i5_not), .in18(i4), .in19(i3), .in20(i2), .in21(i1), .in22(i0_not));
and24$ and_gate186(.out(and186), .in0(i23_not), .in1(i22), .in2(i21
), .in3(i20_not), .in4(i19), .in5(i18), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7_not), .in17(i6), .in18(i5), .in19(i4_not), .in20(i3), .in21(i2), .in22(i1), .in23(i0));
and24$ and_gate187(.out(and187), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15_not), .in9(i14), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1), .in23(i0_not));
and24$ and_gate188(.out(and188), .in0(i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19
), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11), .in13(i10), .in14(i9_not), .in15(i8_not), .in16(i7), .in17(i6), .in18(i5_not), .in19(i4), .in20(i3), .in21(i2), .in22(i1_not), .in23(i0_not));
and21$ and_gate189(.out(and189), .in0(i20_not), .in1(i19), .in2(i18_not), .in3(i17), .in4(i16), .in5(i15_not), .in6(i14), .in7(i13), .in8(i12_not), .in9(i11), .in10(i10), .in11(i9), .in12(i8), .in13(i7_not), .in14(i6_not), .in15(i5), .in16(i4), .in17(i3_not), .in18(i2), .in19(i1), .in20(i0_not));
and21$ and_gate190(.out(and190), .in0(i20_not), .in1(i19), .in2(i18_not), .in3(i17), .in4(i16_not), .in5(i15), .in6(i14), .in7(i13_not), .in8(i12), .in9(i11
), .in10(i10), .in11(i9), .in12(i8), .in13(i7_not), .in14(i6_not), .in15(i5), .in16(i4), .in17(i3_not), .in18(i2_not), .in19(i1), .in20(i0));
and18$ and_gate191(.out(and191), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13_not), .in5(i12_not), .in6(i11_not), .in7(i10_not), .in8(i9), .in9(i8_not), .in10(i7_not), .in11(i6), .in12(i5_not), .in13(i4_not), .in14(i3), .in15(i2), .in16(i1_not), .in17(i0));
and18$ and_gate192(.out(and192), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14
), .in4(i13_not), .in5(i12), .in6(i11_not), .in7(i10_not), .in8(i9), .in9(i8_not), .in10(i7_not), .in11(i6), .in12(i5), .in13(i4_not), .in14(i3), .in15(i2), .in16(i1_not), .in17(i0));
and18$ and_gate193(.out(and193), .in0(i17_not), .in1(i16
), .in2(i15_not), .in3(i14), .in4(i13), .in5(i12_not), .in6(i11), .in7(i10_not), .in8(i9), .in9(i8_not), .in10(i7), .in11(i6), .in12(i5_not), .in13(i4_not), .in14(i3), .in15(i2_not), .in16(i1), .in17(i0));
and18$ and_gate194(.out(and194), .in0(i17_not), .in1(i16), .in2(i15_not), .in3(i14), .in4(i13_not), .in5(i12), .in6(i11), .in7(i10), .in8(i9_not), .in9(i8), .in10(i7), .in11(i6), .in12(i5), .in13(i4_not), .in14(i3_not), .in15(i2), .in16(i1), .in17(i0_not));
and16$ and_gate195(.out(and195), .in0(
i23), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14), .in10(i5_not), .in11(i4), .in12(i3_not), .in13(i2), .in14(i1_not), .in15(i0));
and16$ and_gate196(.out(and196), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19), .in5(i18), .in6(i17_not), .in7(i16_not), .in8(i15), .in9(i14), .in10(i5_not), .in11(i4), .in12(i3_not), .in13(i2), .in14(i1), .in15(i0_not));
and16$ and_gate197(.out(and197), .in0(i23_not), .in1(i22), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18), .in6(i17), .in7(i16_not), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i10), .in14(i9), .in15(i8_not));
and16$ and_gate198(.out(and198), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12_not), .in12(i11_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and16$ and_gate199(.out(and199), .in0(i23_not), .in1(i22_not), .in2(i21), .in3(i20_not), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and16$ and_gate200(.out(and200), .in0(
i23), .in1(i22), .in2(i21), .in3(i20), .in4(i19_not), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15_not), .in9(i14_not), .in10(i13), .in11(i12), .in12(i11_not), .in13(i2_not), .in14(i1), .in15(i0_not));
and16$ and_gate201(.out(and201), .in0(
i23), .in1(i22), .in2(i21_not), .in3(i20_not), .in4(i19), .in5(i18_not), .in6(i17), .in7(i16), .in8(i15), .in9(i14_not), .in10(i5_not), .in11(i4), .in12(i3_not), .in13(i2), .in14(i1_not), .in15(i0_not));
and9$ and_gate202(.out(and202), .in0(i8_not), .in1(i7_not), .in2(i6), .in3(i5), .in4(i4), .in5(i3_not), .in6(i2_not), .in7(i1_not), .in8(i0_not));
and9$ and_gate203(.out(and203), .in0(i8_not), .in1(i7_not), .in2(i6), .in3(i5), .in4(i4_not), .in5(i3), .in6(i2), .in7(i1_not), .in8(i0_not));

or38$ or_gate0(.out(or0), .in0(and0), .in1(and1), .in2(and2), .in3(and3), .in4(and4), .in5(and5), .in6(and6), .in7(and7), .in8(and8), .in9(and9), .in10(and10), .in11(and11), .in12(and12), .in13(and13), .in14(and14), .in15(and15), .in16(and16), .in17(and17), .in18(and18), .in19(and19), .in20(and20), .in21(and21), .in22(and22), .in23(and23), .in24(and24), .in25(and25), .in26(and26), .in27(and27), .in28(and28), .in29(and29), .in30(and30), .in31(and31), .in32(and32), .in33(and33), .in34(and34), .in35(and35), .in36(and36), .in37(and37));
or39$ or_gate1(.out(or1), .in0(and38), .in1(and39), .in2(and40), .in3(and41), .in4(and42), .in5(and43), .in6(and44), .in7(and45), .in8(and46), .in9(and47), .in10(and48), .in11(and49), .in12(and50), .in13(and51), .in14(and52), .in15(and53), .in16(and54), .in17(and55), .in18(and56), .in19(and57), .in20(and58), .in21(and59), .in22(and60), .in23(and61), .in24(and62), .in25(and63), .in26(and64), .in27(and65), .in28(and66), .in29(and67), .in30(and68), .in31(and69), .in32(and70), .in33(and71), .in34(and72), .in35(and73), .in36(and74), .in37(and75), .in38(and76));
or33$ or_gate2(.out(or2), .in0(and77), .in1(and78), .in2(and79), .in3(and80), .in4(and81), .in5(and82), .in6(and83), .in7(and84), .in8(and85), .in9(and86), .in10(and87), .in11(and88), .in12(and89), .in13(and90), .in14(and91), .in15(and92), .in16(and93), .in17(and94), .in18(and95), .in19(and96), .in20(and97), .in21(and98), .in22(and99), .in23(and100), .in24(and101), .in25(and102), .in26(and103), .in27(and104), .in28(and105), .in29(and106), .in30(and107), .in31(and108), .in32(and109));
or32$ or_gate3(.out(or3), .in0(and110), .in1(and111), .in2(and112), .in3(and113), .in4(and114), .in5(and115), .in6(and116), .in7(and117), .in8(and118), .in9(and119), .in10(and120), .in11(and121), .in12(and122), .in13(and123), .in14(and124), .in15(and125), .in16(and126), .in17(and127), .in18(and128), .in19(and129), .in20(and130), .in21(and131), .in22(and132), .in23(and133), .in24(and134), .in25(and135), .in26(and136), .in27(and137), .in28(and138), .in29(and139), .in30(and140), .in31(and141));
or32$ or_gate4(.out(or4), .in0(and142), .in1(and143), .in2(and144), .in3(and145), .in4(and146), .in5(and147), .in6(and148), .in7(and149), .in8(and150), .in9(and151), .in10(and152), .in11(and153), .in12(and154), .in13(and155), .in14(and156), .in15(and157), .in16(and158), .in17(and159), .in18(and160), .in19(and161), .in20(and162), .in21(and163), .in22(and164), .in23(and165), .in24(and166), .in25(and167), .in26(and168), .in27(and169), .in28(and170), .in29(and171), .in30(and172), .in31(and173));
or30$ or_gate5(.out(or5), .in0(and174), .in1(and175), .in2(and176), .in3(and177), .in4(and178), .in5(and179), .in6(and180), .in7(and181), .in8(and182), .in9(and183), .in10(and184), .in11(and185), .in12(and186), .in13(and187), .in14(and188), .in15(and189), .in16(and190), .in17(and191), .in18(and192), .in19(and193), .in20(and194), .in21(and195), .in22(and196), .in23(and197), .in24(and198), .in25(and199), .in26(and200), .in27(and201), .in28(and202), .in29(and203));

assign pre_seg_override_valid = or0;
assign pre_seg_override[2] = or1;
assign pre_seg_override[1] = or2;
assign pre_seg_override[0] = or3;
assign pre_repeat = or4;
assign pre_size_override = or5;


endmodule
   
