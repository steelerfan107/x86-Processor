module opcode_modrm_control_cloud (
input modrm7, 
input modrm6, 
input modrm5, 
input modrm4, 
input modrm3, 
input modrm2, 
input modrm1, 
input modrm0, 
input op15, 
input op14, 
input op13, 
input op12, 
input op11, 
input op10, 
input op9, 
input op8, 
input op7, 
input op6, 
input op5, 
input op4, 
input op3, 
input op2, 
input op1, 
input op0,
output setd, 
output cleard, 
output size2, 
output size1, 
output size0, 
output op0_2, 
output op0_1, 
output op0_0, 
output op1_2, 
output op1_1, 
output op1_0, 
output op0_reg_4, 
output op0_reg_3, 
output op0_reg_2, 
output op0_reg_1, 
output op0_reg_0, 
output op1_reg_4, 
output op1_reg_3, 
output op1_reg_2, 
output op1_reg_1, 
output op1_reg_0, 
output alu_op_3, 
output alu_op_2, 
output alu_op_1, 
output alu_op_0, 
output flag0_2, 
output flag0_1, 
output flag0_0, 
output flag1_2, 
output flag1_1, 
output flag1_0, 
output stack_op_1, 
output stack_op_0, 
output rom_control_2, 
output rom_control_1, 
output rom_control_0				   
);

wire modrm7_not;
wire modrm6_not;
wire modrm5_not;
wire modrm4_not;
wire modrm3_not;
wire op13_not;
wire op12_not;
wire op11_not;
wire op10_not;
wire op9_not;
wire and0;
wire op15_not;
wire op14_not;
wire op8_not;
wire op6_not;
wire op5_not;
wire op2_not;
wire op0_not;
wire and1;
wire modrm2_not;
wire modrm1_not;
wire modrm0_not;
wire and2;
wire op12_not;
wire op7_not;
wire op4_not;
wire and3;
wire op14_not;
wire op1_not;
wire and4;
wire op15_not;
wire and5;
wire and6;
wire or0;
wire and7;
wire modrm5_not;
wire modrm0_not;
wire and8;
wire and9;
wire modrm6_not;
wire and10;
wire modrm2_not;
wire and11;
wire modrm7_not;
wire and12;
wire modrm4_not;
wire and13;
wire and14;
wire and15;
wire and16;
wire op13_not;
wire op3_not;
wire and17;
wire modrm7_not;
wire and18;
wire op11_not;
wire and19;
wire op8_not;
wire and20;
wire and21;
wire and22;
wire and23;
wire op15_not;
wire op2_not;
wire and24;
wire op5_not;
wire and25;
wire op9_not;
wire and26;
wire and27;
wire op6_not;
wire and28;
wire op10_not;
wire and29;
wire and30;
wire and31;
wire and32;
wire and33;
wire and34;
wire and35;
wire op7_not;
wire and36;
wire and37;
wire and38;
wire and39;
wire and40;
wire and41;
wire and42;
wire and43;
wire and44;
wire or1;
wire and45;
wire and46;
wire and47;
wire op1_not;
wire and48;
wire modrm1_not;
wire and49;
wire and50;
wire and51;
wire and52;
wire and53;
wire and54;
wire and55;
wire and56;
wire and57;
wire and58;
wire and59;
wire and60;
wire op3_not;
wire and61;
wire and62;
wire and63;
wire and64;
wire and65;
wire and66;
wire and67;
wire and68;
wire and69;
wire and70;
wire and71;
wire and72;
wire and73;
wire and74;
wire and75;
wire or2;
wire and76;
wire and77;
wire and78;
wire and79;
wire and80;
wire and81;
wire and82;
wire and83;
wire and84;
wire and85;
wire and86;
wire and87;
wire and88;
wire and89;
wire modrm3_not;
wire and90;
wire and91;
wire and92;
wire and93;
wire and94;
wire and95;
wire and96;
wire and97;
wire and98;
wire and99;
wire and100;
wire and101;
wire and102;
wire and103;
wire and104;
wire op4_not;
wire and105;
wire and106;
wire and107;
wire and108;
wire and109;
wire and110;
wire or3;
wire and111;
wire and112;
wire and113;
wire and114;
wire and115;
wire and116;
wire and117;
wire and118;
wire and119;
wire and120;
wire and121;
wire and122;
wire or4;
wire and123;
wire and124;
wire and125;
wire and126;
wire and127;
wire and128;
wire and129;
wire and130;
wire and131;
wire and132;
wire and133;
wire and134;
wire and135;
wire and136;
wire and137;
wire and138;
wire and139;
wire and140;
wire and141;
wire and142;
wire and143;
wire and144;
wire and145;
wire and146;
wire and147;
wire and148;
wire or5;
wire and149;
wire and150;
wire and151;
wire and152;
wire and153;
wire and154;
wire and155;
wire and156;
wire and157;
wire and158;
wire and159;
wire and160;
wire and161;
wire and162;
wire and163;
wire and164;
wire and165;
wire and166;
wire and167;
wire and168;
wire and169;
wire and170;
wire and171;
wire and172;
wire and173;
wire and174;
wire and175;
wire and176;
wire and177;
wire and178;
wire and179;
wire or6;
wire and180;
wire and181;
wire or7;
wire and182;
wire and183;
wire and184;
wire and185;
wire and186;
wire and187;
wire and188;
wire and189;
wire and190;
wire and191;
wire and192;
wire and193;
wire and194;
wire and195;
wire and196;
wire and197;
wire and198;
wire and199;
wire and200;
wire and201;
wire and202;
wire and203;
wire and204;
wire and205;
wire and206;
wire and207;
wire and208;
wire and209;
wire and210;
wire or8;
wire and211;
wire and212;
wire and213;
wire and214;
wire and215;
wire and216;
wire and217;
wire and218;
wire and219;
wire and220;
wire and221;
wire and222;
wire and223;
wire and224;
wire or9;
wire and225;
wire and226;
wire and227;
wire and228;
wire or10;
wire and229;
wire and230;
wire and231;
wire or11;
wire and232;
wire and233;
wire and234;
wire and235;
wire or12;
wire and236;
wire and237;
wire and238;
wire and239;
wire and240;
wire and241;
wire and242;
wire and243;
wire and244;
wire and245;
wire and246;
wire and247;
wire or13;
wire and248;
wire and249;
wire or14;
wire and250;
wire and251;
wire and252;
wire and253;
wire and254;
wire and255;
wire and256;
wire and257;
wire and258;
wire and259;
wire and260;
wire and261;
wire and262;
wire and263;
wire and264;
wire and265;
wire and266;
wire or15;
wire and267;
wire and268;
wire and269;
wire and270;
wire and271;
wire and272;
wire and273;
wire and274;
wire and275;
wire and276;
wire and277;
wire and278;
wire and279;
wire and280;
wire and281;
wire and282;
wire and283;
wire and284;
wire and285;
wire and286;
wire and287;
wire and288;
wire and289;
wire and290;
wire or16;
wire and291;
wire and292;
wire and293;
wire and294;
wire and295;
wire and296;
wire and297;
wire and298;
wire and299;
wire and300;
wire and301;
wire and302;
wire and303;
wire and304;
wire and305;
wire and306;
wire and307;
wire and308;
wire and309;
wire and310;
wire and311;
wire or17;
wire and312;
wire and313;
wire and314;
wire and315;
wire and316;
wire and317;
wire and318;
wire and319;
wire and320;
wire and321;
wire and322;
wire and323;
wire or18;
wire and324;
wire and325;
wire and326;
wire and327;
wire and328;
wire and329;
wire or19;
wire and330;
wire and331;
wire and332;
wire and333;
wire and334;
wire or20;
wire and335;
wire and336;
wire or21;
wire and337;
wire and338;
wire and339;
wire and340;
wire and341;
wire and342;
wire and343;
wire and344;
wire or22;
wire and345;
wire and346;
wire and347;
wire and348;
wire and349;
wire and350;
wire and351;
wire or23;
wire and352;
wire and353;
wire and354;
wire or24;
wire and355;
wire and356;
wire and357;
wire or25;
wire and358;
wire and359;
wire and360;
wire and361;
wire and362;
wire or26;

inv1$ modrm7_inv (.out(modrm7_not), .in(modrm7));
inv1$ modrm6_inv (.out(modrm6_not), .in(modrm6));
inv1$ modrm5_inv (.out(modrm5_not), .in(modrm5));
inv1$ modrm4_inv (.out(modrm4_not), .in(modrm4));
inv1$ modrm3_inv (.out(modrm3_not), .in(modrm3));
inv1$ op13_inv (.out(op13_not), .in(op13));
inv1$ op12_inv (.out(op12_not), .in(op12));
inv1$ op11_inv (.out(op11_not), .in(op11));
inv1$ op10_inv (.out(op10_not), .in(op10));
inv1$ op9_inv (.out(op9_not), .in(op9));
inv1$ op15_inv (.out(op15_not), .in(op15));
inv1$ op14_inv (.out(op14_not), .in(op14));
inv1$ op8_inv (.out(op8_not), .in(op8));
inv1$ op6_inv (.out(op6_not), .in(op6));
inv1$ op5_inv (.out(op5_not), .in(op5));
inv1$ op2_inv (.out(op2_not), .in(op2));
inv1$ op0_inv (.out(op0_not), .in(op0));
inv1$ modrm2_inv (.out(modrm2_not), .in(modrm2));
inv1$ modrm1_inv (.out(modrm1_not), .in(modrm1));
inv1$ modrm0_inv (.out(modrm0_not), .in(modrm0));
inv1$ op12_inv (.out(op12_not), .in(op12));
inv1$ op7_inv (.out(op7_not), .in(op7));
inv1$ op4_inv (.out(op4_not), .in(op4));
inv1$ op14_inv (.out(op14_not), .in(op14));
inv1$ op1_inv (.out(op1_not), .in(op1));
inv1$ op15_inv (.out(op15_not), .in(op15));
inv1$ modrm5_inv (.out(modrm5_not), .in(modrm5));
inv1$ modrm0_inv (.out(modrm0_not), .in(modrm0));
inv1$ modrm6_inv (.out(modrm6_not), .in(modrm6));
inv1$ modrm2_inv (.out(modrm2_not), .in(modrm2));
inv1$ modrm7_inv (.out(modrm7_not), .in(modrm7));
inv1$ modrm4_inv (.out(modrm4_not), .in(modrm4));
inv1$ op13_inv (.out(op13_not), .in(op13));
inv1$ op3_inv (.out(op3_not), .in(op3));
inv1$ modrm7_inv (.out(modrm7_not), .in(modrm7));
inv1$ op11_inv (.out(op11_not), .in(op11));
inv1$ op8_inv (.out(op8_not), .in(op8));
inv1$ op15_inv (.out(op15_not), .in(op15));
inv1$ op2_inv (.out(op2_not), .in(op2));
inv1$ op5_inv (.out(op5_not), .in(op5));
inv1$ op9_inv (.out(op9_not), .in(op9));
inv1$ op6_inv (.out(op6_not), .in(op6));
inv1$ op10_inv (.out(op10_not), .in(op10));
inv1$ op7_inv (.out(op7_not), .in(op7));
inv1$ op1_inv (.out(op1_not), .in(op1));
inv1$ modrm1_inv (.out(modrm1_not), .in(modrm1));
inv1$ op3_inv (.out(op3_not), .in(op3));
inv1$ modrm3_inv (.out(modrm3_not), .in(modrm3));
inv1$ op4_inv (.out(op4_not), .in(op4));

and16$ and_gate0(.out(and0), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0), .in8(op15
), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8));
and16$ and_gate1(.out(and1), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4
), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate2(.out(and2), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate3(.out(and3), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate4(.out(and4), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and15$ and_gate5(.out(and5), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op3), .in12(op2), .in13(op1), .in14(op0_not));
and16$ and_gate6(.out(and6), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3
), .in13(op2_not), .in14(op1), .in15(op0));
and16$ and_gate7(.out(and7), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate8(.out(and8), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11), .in13(op10
), .in14(op9), .in15(op8));
and16$ and_gate9(.out(and9), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1
), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8_not));
and15$ and_gate10(.out(and10), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12
), .in12(op11_not), .in13(op10_not), .in14(op8));
and16$ and_gate11(.out(and11), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11), .in13(op10), .in14(op9), .in15(op8));
and15$ and_gate12(.out(and12), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14
), .in10(op13_not), .in11(op12), .in12(op11_not), .in13(op10_not), .in14(op8));
and16$ and_gate13(.out(and13), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10), .in14(op9
), .in15(op8_not));
and16$ and_gate14(.out(and14), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4
), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate15(.out(and15), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7
), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate16(.out(and16), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10
), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1_not), .in15(op0));
and16$ and_gate17(.out(and17), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate18(.out(and18), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0), .in8(op15
), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8_not));
and16$ and_gate19(.out(and19), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8_not));
and16$ and_gate20(.out(and20), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate21(.out(and21), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11
), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and15$ and_gate22(.out(and22), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and15$ and_gate23(.out(and23), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and16$ and_gate24(.out(and24), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate25(.out(and25), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate26(.out(and26), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0));
and15$ and_gate27(.out(and27), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and16$ and_gate28(.out(and28), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0_not));
and15$ and_gate29(.out(and29), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1_not));
and16$ and_gate30(.out(and30), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate31(.out(and31), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate32(.out(and32), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6
), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate33(.out(and33), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate34(.out(and34), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate35(.out(and35), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3
), .in13(op2_not), .in14(op1), .in15(op0));
and16$ and_gate36(.out(and36), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate37(.out(and37), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and15$ and_gate38(.out(and38), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op0));
and15$ and_gate39(.out(and39), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate40(.out(and40), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate41(.out(and41), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1), .in14(op0_not));
and15$ and_gate42(.out(and42), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not), .in14(op0_not));
and15$ and_gate43(.out(and43), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1));
and15$ and_gate44(.out(and44), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1));
and16$ and_gate45(.out(and45), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate46(.out(and46), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate47(.out(and47), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate48(.out(and48), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate49(.out(and49), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and16$ and_gate50(.out(and50), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and16$ and_gate51(.out(and51), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9
), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate52(.out(and52), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and14$ and_gate53(.out(and53), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2
), .in6(modrm1), .in7(modrm0), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12), .in12(op11_not), .in13(op10_not));
and14$ and_gate54(.out(and54), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12
), .in12(op11_not), .in13(op10_not));
and16$ and_gate55(.out(and55), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2
), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8));
and16$ and_gate56(.out(and56), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1
), .in15(op0));
and16$ and_gate57(.out(and57), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op4
), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate58(.out(and58), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate59(.out(and59), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate60(.out(and60), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate61(.out(and61), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and15$ and_gate62(.out(and62), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6
), .in10(op5), .in11(op3), .in12(op2), .in13(op1), .in14(op0_not));
and16$ and_gate63(.out(and63), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate64(.out(and64), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0));
and16$ and_gate65(.out(and65), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2
), .in14(op1), .in15(op0_not));
and16$ and_gate66(.out(and66), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6
), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate67(.out(and67), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate68(.out(and68), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0));
and15$ and_gate69(.out(and69), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1), .in14(op0_not));
and15$ and_gate70(.out(and70), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0));
and15$ and_gate71(.out(and71), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1_not), .in14(op0));
and15$ and_gate72(.out(and72), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not), .in14(op0));
and5$ and_gate73(.out(and73), .in0(op15_not), .in1(op14), .in2(op13_not), .in3(op12), .in4(op11));
and5$ and_gate74(.out(and74), .in0(op15), .in1(op14_not), .in2(op13), .in3(op12), .in4(op11));
and5$ and_gate75(.out(and75), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and16$ and_gate76(.out(and76), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8_not));
and16$ and_gate77(.out(and77), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8_not));
and16$ and_gate78(.out(and78), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and16$ and_gate79(.out(and79), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15
), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and16$ and_gate80(.out(and80), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate81(.out(and81), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate82(.out(and82), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15
), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and16$ and_gate83(.out(and83), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1_not), .in15(op0));
and14$ and_gate84(.out(and84), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12), .in12(op11_not), .in13(op10_not));
and14$ and_gate85(.out(and85), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2
), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12), .in12(op11_not), .in13(op10_not));
and16$ and_gate86(.out(and86), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8));
and16$ and_gate87(.out(and87), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8
), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate88(.out(and88), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11
), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate89(.out(and89), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8_not));
and16$ and_gate90(.out(and90), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8_not));
and16$ and_gate91(.out(and91), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate92(.out(and92), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and15$ and_gate93(.out(and93), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and15$ and_gate94(.out(and94), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15
), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and16$ and_gate95(.out(and95), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11
), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and15$ and_gate96(.out(and96), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and15$ and_gate97(.out(and97), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1_not));
and16$ and_gate98(.out(and98), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate99(.out(and99), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate100(.out(and100), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3
), .in13(op2_not), .in14(op1), .in15(op0));
and16$ and_gate101(.out(and101), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7
), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate102(.out(and102), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and15$ and_gate103(.out(and103), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1), .in14(op0_not));
and15$ and_gate104(.out(and104), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op0));
and15$ and_gate105(.out(and105), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate106(.out(and106), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate107(.out(and107), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not), .in14(op0));
and15$ and_gate108(.out(and108), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1));
and5$ and_gate109(.out(and109), .in0(
op15), .in1(op14_not), .in2(op13), .in3(op12), .in4(op11));
and5$ and_gate110(.out(and110), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and16$ and_gate111(.out(and111), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate112(.out(and112), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate113(.out(and113), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and16$ and_gate114(.out(and114), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4
), .in12(op3), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate115(.out(and115), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7
), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate116(.out(and116), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate117(.out(and117), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and15$ and_gate118(.out(and118), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op3), .in12(op2), .in13(op1), .in14(op0_not));
and15$ and_gate119(.out(and119), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4), .in12(op2
), .in13(op1), .in14(op0));
and14$ and_gate120(.out(and120), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op2), .in12(op1), .in13(op0_not));
and16$ and_gate121(.out(and121), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0));
and5$ and_gate122(.out(and122), .in0(op15_not), .in1(op14), .in2(op13_not), .in3(op12), .in4(op11));
and16$ and_gate123(.out(and123), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate124(.out(and124), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate125(.out(and125), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate126(.out(and126), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14
), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate127(.out(and127), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10
), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and16$ and_gate128(.out(and128), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate129(.out(and129), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0));
and16$ and_gate130(.out(and130), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate131(.out(and131), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8
), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and15$ and_gate132(.out(and132), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op3), .in12(op2), .in13(op1), .in14(op0_not));
and16$ and_gate133(.out(and133), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate134(.out(and134), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate135(.out(and135), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate136(.out(and136), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate137(.out(and137), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate138(.out(and138), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate139(.out(and139), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0));
and16$ and_gate140(.out(and140), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1), .in15(op0_not));
and16$ and_gate141(.out(and141), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate142(.out(and142), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3
), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate143(.out(and143), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0));
and15$ and_gate144(.out(and144), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0));
and15$ and_gate145(.out(and145), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1_not), .in14(op0));
and15$ and_gate146(.out(and146), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1), .in14(op0_not));
and15$ and_gate147(.out(and147), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not), .in14(op0_not));
and15$ and_gate148(.out(and148), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1));
and16$ and_gate149(.out(and149), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8));
and15$ and_gate150(.out(and150), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12), .in12(op11_not), .in13(op10_not), .in14(op9));
and15$ and_gate151(.out(and151), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12), .in12(op11_not), .in13(op10_not), .in14(op9));
and16$ and_gate152(.out(and152), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate153(.out(and153), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8_not));
and16$ and_gate154(.out(and154), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2
), .in14(op1), .in15(op0));
and16$ and_gate155(.out(and155), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8));
and16$ and_gate156(.out(and156), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate157(.out(and157), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0), .in8(op15
), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8_not));
and16$ and_gate158(.out(and158), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8_not));
and15$ and_gate159(.out(and159), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and15$ and_gate160(.out(and160), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and15$ and_gate161(.out(and161), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and15$ and_gate162(.out(and162), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op3
), .in12(op2), .in13(op1), .in14(op0_not));
and16$ and_gate163(.out(and163), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7
), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate164(.out(and164), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate165(.out(and165), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate166(.out(and166), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0));
and16$ and_gate167(.out(and167), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate168(.out(and168), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0));
and16$ and_gate169(.out(and169), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3
), .in13(op2), .in14(op1), .in15(op0_not));
and16$ and_gate170(.out(and170), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate171(.out(and171), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate172(.out(and172), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1
), .in15(op0));
and15$ and_gate173(.out(and173), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0));
and15$ and_gate174(.out(and174), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1_not), .in14(op0));
and15$ and_gate175(.out(and175), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1), .in14(op0_not));
and15$ and_gate176(.out(and176), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not), .in14(op0_not));
and15$ and_gate177(.out(and177), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2
), .in13(op1_not), .in14(op0));
and15$ and_gate178(.out(and178), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1));
and5$ and_gate179(.out(and179), .in0(op15), .in1(op14_not), .in2(op13), .in3(op12), .in4(op11));
and16$ and_gate180(.out(and180), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3
), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate181(.out(and181), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6
), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate182(.out(and182), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate183(.out(and183), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8_not));
and16$ and_gate184(.out(and184), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and16$ and_gate185(.out(and185), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15
), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and16$ and_gate186(.out(and186), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and14$ and_gate187(.out(and187), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2
), .in6(modrm1), .in7(modrm0), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12), .in12(op11_not), .in13(op10_not));
and14$ and_gate188(.out(and188), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12
), .in12(op11_not), .in13(op10_not));
and16$ and_gate189(.out(and189), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2
), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8));
and16$ and_gate190(.out(and190), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1
), .in15(op0));
and16$ and_gate191(.out(and191), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4
), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate192(.out(and192), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8_not));
and16$ and_gate193(.out(and193), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15
), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8_not));
and16$ and_gate194(.out(and194), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and15$ and_gate195(.out(and195), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and15$ and_gate196(.out(and196), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and15$ and_gate197(.out(and197), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and16$ and_gate198(.out(and198), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate199(.out(and199), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3
), .in13(op2), .in14(op1), .in15(op0_not));
and16$ and_gate200(.out(and200), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate201(.out(and201), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate202(.out(and202), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1
), .in15(op0));
and15$ and_gate203(.out(and203), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1), .in14(op0_not));
and15$ and_gate204(.out(and204), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate205(.out(and205), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate206(.out(and206), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not), .in14(op0_not));
and15$ and_gate207(.out(and207), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2
), .in13(op1_not), .in14(op0));
and15$ and_gate208(.out(and208), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1));
and5$ and_gate209(.out(and209), .in0(op15), .in1(op14_not), .in2(op13), .in3(op12), .in4(op11));
and5$ and_gate210(.out(and210), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and16$ and_gate211(.out(and211), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate212(.out(and212), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate213(.out(and213), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate214(.out(and214), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6
), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and15$ and_gate215(.out(and215), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9
), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op3), .in12(op2), .in13(op1), .in14(op0_not));
and16$ and_gate216(.out(and216), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate217(.out(and217), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate218(.out(and218), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate219(.out(and219), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0));
and16$ and_gate220(.out(and220), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1), .in15(op0_not));
and15$ and_gate221(.out(and221), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0));
and15$ and_gate222(.out(and222), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1_not), .in14(op0));
and15$ and_gate223(.out(and223), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1), .in14(op0_not));
and15$ and_gate224(.out(and224), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1));
and16$ and_gate225(.out(and225), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate226(.out(and226), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8
), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and16$ and_gate227(.out(and227), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and15$ and_gate228(.out(and228), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1
), .in14(op0_not));
and16$ and_gate229(.out(and229), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0_not));
and14$ and_gate230(.out(and230), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op1), .in13(op0_not));
and16$ and_gate231(.out(and231), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate232(.out(and232), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate233(.out(and233), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8
), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and16$ and_gate234(.out(and234), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0_not));
and16$ and_gate235(.out(and235), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate236(.out(and236), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5
), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate237(.out(and237), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and16$ and_gate238(.out(and238), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and16$ and_gate239(.out(and239), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and16$ and_gate240(.out(and240), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2
), .in14(op1), .in15(op0));
and16$ and_gate241(.out(and241), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5
), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate242(.out(and242), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9
), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and15$ and_gate243(.out(and243), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1), .in14(op0_not));
and15$ and_gate244(.out(and244), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate245(.out(and245), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate246(.out(and246), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1));
and5$ and_gate247(.out(and247), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and14$ and_gate248(.out(and248), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0
), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12), .in12(op11_not), .in13(op10_not));
and14$ and_gate249(.out(and249), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12), .in12(op11_not), .in13(op10_not));
and16$ and_gate250(.out(and250), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate251(.out(and251), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and14$ and_gate252(.out(and252), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2
), .in6(modrm1), .in7(modrm0), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12), .in12(op11_not), .in13(op10_not));
and14$ and_gate253(.out(and253), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12
), .in12(op11_not), .in13(op10_not));
and16$ and_gate254(.out(and254), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2
), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8));
and16$ and_gate255(.out(and255), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate256(.out(and256), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0), .in8(op15
), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8_not));
and16$ and_gate257(.out(and257), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8_not));
and15$ and_gate258(.out(and258), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and15$ and_gate259(.out(and259), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op3), .in12(op2), .in13(op1), .in14(op0_not));
and16$ and_gate260(.out(and260), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3
), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate261(.out(and261), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7
), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and14$ and_gate262(.out(and262), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2_not));
and16$ and_gate263(.out(and263), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate264(.out(and264), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3
), .in13(op2), .in14(op1_not), .in15(op0));
and15$ and_gate265(.out(and265), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7
), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1));
and5$ and_gate266(.out(and266), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and16$ and_gate267(.out(and267), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate268(.out(and268), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8_not));
and16$ and_gate269(.out(and269), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and14$ and_gate270(.out(and270), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12), .in12(op11_not), .in13(op10_not));
and14$ and_gate271(.out(and271), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15
), .in9(op14), .in10(op13_not), .in11(op12), .in12(op11_not), .in13(op10_not));
and16$ and_gate272(.out(and272), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8));
and16$ and_gate273(.out(and273), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4
), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate274(.out(and274), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8_not));
and16$ and_gate275(.out(and275), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15
), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8_not));
and16$ and_gate276(.out(and276), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate277(.out(and277), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1
), .in15(op0));
and16$ and_gate278(.out(and278), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate279(.out(and279), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate280(.out(and280), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate281(.out(and281), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate282(.out(and282), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate283(.out(and283), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and15$ and_gate284(.out(and284), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op2_not), .in13(op1), .in14(op0));
and16$ and_gate285(.out(and285), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate286(.out(and286), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate287(.out(and287), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1), .in15(op0));
and15$ and_gate288(.out(and288), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op0));
and15$ and_gate289(.out(and289), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1));
and5$ and_gate290(.out(and290), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and16$ and_gate291(.out(and291), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate292(.out(and292), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8_not));
and16$ and_gate293(.out(and293), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2
), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and16$ and_gate294(.out(and294), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate295(.out(and295), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2
), .in14(op1), .in15(op0));
and16$ and_gate296(.out(and296), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and15$ and_gate297(.out(and297), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and16$ and_gate298(.out(and298), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and15$ and_gate299(.out(and299), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6
), .in10(op5), .in11(op3), .in12(op2), .in13(op1), .in14(op0_not));
and16$ and_gate300(.out(and300), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate301(.out(and301), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and15$ and_gate302(.out(and302), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op2_not), .in13(op1
), .in14(op0));
and16$ and_gate303(.out(and303), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5
), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate304(.out(and304), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0));
and14$ and_gate305(.out(and305), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op1_not));
and16$ and_gate306(.out(and306), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate307(.out(and307), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0));
and15$ and_gate308(.out(and308), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7
), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op0));
and15$ and_gate309(.out(and309), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1));
and15$ and_gate310(.out(and310), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1));
and5$ and_gate311(.out(and311), .in0(
op15), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and16$ and_gate312(.out(and312), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11_not), .in13(op10), .in14(op9), .in15(op8_not));
and16$ and_gate313(.out(and313), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and16$ and_gate314(.out(and314), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9), .in15(op8));
and14$ and_gate315(.out(and315), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12), .in12(op11_not), .in13(op10_not));
and16$ and_gate316(.out(and316), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15
), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8));
and16$ and_gate317(.out(and317), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1), .in7(modrm0), .in8(op15), .in9(op14), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not), .in15(op8_not));
and16$ and_gate318(.out(and318), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0));
and15$ and_gate319(.out(and319), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11_not), .in13(op10_not), .in14(op9_not));
and15$ and_gate320(.out(and320), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5
), .in11(op3), .in12(op2), .in13(op1), .in14(op0_not));
and16$ and_gate321(.out(and321), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and14$ and_gate322(.out(and322), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op1_not));
and16$ and_gate323(.out(and323), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1
), .in15(op0));
and16$ and_gate324(.out(and324), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate325(.out(and325), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate326(.out(and326), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11
), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate327(.out(and327), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate328(.out(and328), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate329(.out(and329), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7
), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate330(.out(and330), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate331(.out(and331), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate332(.out(and332), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate333(.out(and333), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate334(.out(and334), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3
), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate335(.out(and335), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4
), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate336(.out(and336), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate337(.out(and337), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(modrm1_not), .in7(modrm0_not), .in8(op15), .in9(op14_not), .in10(op13_not), .in11(op12_not), .in12(op11), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate338(.out(and338), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and16$ and_gate339(.out(and339), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0_not));
and16$ and_gate340(.out(and340), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate341(.out(and341), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0));
and15$ and_gate342(.out(and342), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4), .in12(op2), .in13(op1), .in14(op0));
and16$ and_gate343(.out(and343), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and5$ and_gate344(.out(and344), .in0(op15_not), .in1(op14), .in2(op13_not), .in3(op12), .in4(op11));
and16$ and_gate345(.out(and345), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(modrm1
), .in7(modrm0_not), .in8(op15), .in9(op14), .in10(op13), .in11(op12), .in12(op11), .in13(op10), .in14(op9), .in15(op8));
and16$ and_gate346(.out(and346), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate347(.out(and347), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1_not), .in15(op0));
and16$ and_gate348(.out(and348), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6
), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate349(.out(and349), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0_not));
and14$ and_gate350(.out(and350), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op2), .in12(op1), .in13(op0_not));
and5$ and_gate351(.out(and351), .in0(op15_not), .in1(op14), .in2(op13_not), .in3(op12), .in4(op11));
and16$ and_gate352(.out(and352), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0));
and16$ and_gate353(.out(and353), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));
and15$ and_gate354(.out(and354), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op2_not), .in13(op1), .in14(op0));
and16$ and_gate355(.out(and355), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5
), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate356(.out(and356), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate357(.out(and357), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate358(.out(and358), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5
), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate359(.out(and359), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2), .in14(op1), .in15(op0));
and16$ and_gate360(.out(and360), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6), .in10(op5_not), .in11(op4_not), .in12(op3), .in13(op2_not), .in14(op1), .in15(op0));
and16$ and_gate361(.out(and361), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4_not), .in12(op3_not), .in13(op2
), .in14(op1_not), .in15(op0_not));
and16$ and_gate362(.out(and362), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6
), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1), .in15(op0_not));

or5$ or_gate0(.out(or0), .in0(and2), .in1(and3), .in2(and4), .in3(and5), .in4(and6));
or38$ or_gate1(.out(or1), .in0(and7), .in1(and8), .in2(and9), .in3(and10), .in4(and11), .in5(and12), .in6(and13), .in7(and14), .in8(and15), .in9(and16), .in10(and17), .in11(and18), .in12(and19), .in13(and20), .in14(and21), .in15(and22), .in16(and23), .in17(and24), .in18(and25), .in19(and26), .in20(and27), .in21(and28), .in22(and29), .in23(and30), .in24(and31), .in25(and32), .in26(and33), .in27(and34), .in28(and35), .in29(and36), .in30(and37), .in31(and38), .in32(and39), .in33(and40), .in34(and41), .in35(and42), .in36(and43), .in37(and44));
or31$ or_gate2(.out(or2), .in0(and45), .in1(and46), .in2(and47), .in3(and48), .in4(and49), .in5(and50), .in6(and51), .in7(and52), .in8(and53), .in9(and54), .in10(and55), .in11(and56), .in12(and57), .in13(and58), .in14(and59), .in15(and60), .in16(and61), .in17(and62), .in18(and63), .in19(and64), .in20(and65), .in21(and66), .in22(and67), .in23(and68), .in24(and69), .in25(and70), .in26(and71), .in27(and72), .in28(and73), .in29(and74), .in30(and75));
or35$ or_gate3(.out(or3), .in0(and76), .in1(and77), .in2(and78), .in3(and79), .in4(and80), .in5(and81), .in6(and82), .in7(and83), .in8(and84), .in9(and85), .in10(and86), .in11(and87), .in12(and88), .in13(and89), .in14(and90), .in15(and91), .in16(and92), .in17(and93), .in18(and94), .in19(and95), .in20(and96), .in21(and97), .in22(and98), .in23(and99), .in24(and100), .in25(and101), .in26(and102), .in27(and103), .in28(and104), .in29(and105), .in30(and106), .in31(and107), .in32(and108), .in33(and109), .in34(and110));
or12$ or_gate4(.out(or4), .in0(and111), .in1(and112), .in2(and113), .in3(and114), .in4(and115), .in5(and116), .in6(and117), .in7(and118), .in8(and119), .in9(and120), .in10(and121), .in11(and122));
or26$ or_gate5(.out(or5), .in0(and123), .in1(and124), .in2(and125), .in3(and126), .in4(and127), .in5(and128), .in6(and129), .in7(and130), .in8(and131), .in9(and132), .in10(and133), .in11(and134), .in12(and135), .in13(and136), .in14(and137), .in15(and138), .in16(and139), .in17(and140), .in18(and141), .in19(and142), .in20(and143), .in21(and144), .in22(and145), .in23(and146), .in24(and147), .in25(and148));
or31$ or_gate6(.out(or6), .in0(and149), .in1(and150), .in2(and151), .in3(and152), .in4(and153), .in5(and154), .in6(and155), .in7(and156), .in8(and157), .in9(and158), .in10(and159), .in11(and160), .in12(and161), .in13(and162), .in14(and163), .in15(and164), .in16(and165), .in17(and166), .in18(and167), .in19(and168), .in20(and169), .in21(and170), .in22(and171), .in23(and172), .in24(and173), .in25(and174), .in26(and175), .in27(and176), .in28(and177), .in29(and178), .in30(and179));
or2$ or_gate7(.out(or7), .in0(and180), .in1(and181));
or29$ or_gate8(.out(or8), .in0(and182), .in1(and183), .in2(and184), .in3(and185), .in4(and186), .in5(and187), .in6(and188), .in7(and189), .in8(and190), .in9(and191), .in10(and192), .in11(and193), .in12(and194), .in13(and195), .in14(and196), .in15(and197), .in16(and198), .in17(and199), .in18(and200), .in19(and201), .in20(and202), .in21(and203), .in22(and204), .in23(and205), .in24(and206), .in25(and207), .in26(and208), .in27(and209), .in28(and210));
or13$ or_gate9(.out(or9), .in0(and212), .in1(and213), .in2(and214), .in3(and215), .in4(and216), .in5(and217), .in6(and218), .in7(and219), .in8(and220), .in9(and221), .in10(and222), .in11(and223), .in12(and224));
or4$ or_gate10(.out(or10), .in0(and225), .in1(and226), .in2(and227), .in3(and228));
or3$ or_gate11(.out(or11), .in0(and229), .in1(and230), .in2(and231));
or4$ or_gate12(.out(or12), .in0(and232), .in1(and233), .in2(and234), .in3(and235));
or11$ or_gate13(.out(or13), .in0(and237), .in1(and238), .in2(and239), .in3(and240), .in4(and241), .in5(and242), .in6(and243), .in7(and244), .in8(and245), .in9(and246), .in10(and247));
or2$ or_gate14(.out(or14), .in0(and248), .in1(and249));
or17$ or_gate15(.out(or15), .in0(and250), .in1(and251), .in2(and252), .in3(and253), .in4(and254), .in5(and255), .in6(and256), .in7(and257), .in8(and258), .in9(and259), .in10(and260), .in11(and261), .in12(and262), .in13(and263), .in14(and264), .in15(and265), .in16(and266));
or24$ or_gate16(.out(or16), .in0(and267), .in1(and268), .in2(and269), .in3(and270), .in4(and271), .in5(and272), .in6(and273), .in7(and274), .in8(and275), .in9(and276), .in10(and277), .in11(and278), .in12(and279), .in13(and280), .in14(and281), .in15(and282), .in16(and283), .in17(and284), .in18(and285), .in19(and286), .in20(and287), .in21(and288), .in22(and289), .in23(and290));
or21$ or_gate17(.out(or17), .in0(and291), .in1(and292), .in2(and293), .in3(and294), .in4(and295), .in5(and296), .in6(and297), .in7(and298), .in8(and299), .in9(and300), .in10(and301), .in11(and302), .in12(and303), .in13(and304), .in14(and305), .in15(and306), .in16(and307), .in17(and308), .in18(and309), .in19(and310), .in20(and311));
or12$ or_gate18(.out(or18), .in0(and312), .in1(and313), .in2(and314), .in3(and315), .in4(and316), .in5(and317), .in6(and318), .in7(and319), .in8(and320), .in9(and321), .in10(and322), .in11(and323));
or6$ or_gate19(.out(or19), .in0(and324), .in1(and325), .in2(and326), .in3(and327), .in4(and328), .in5(and329));
or5$ or_gate20(.out(or20), .in0(and330), .in1(and331), .in2(and332), .in3(and333), .in4(and334));
or2$ or_gate21(.out(or21), .in0(and335), .in1(and336));
or8$ or_gate22(.out(or22), .in0(and337), .in1(and338), .in2(and339), .in3(and340), .in4(and341), .in5(and342), .in6(and343), .in7(and344));
or7$ or_gate23(.out(or23), .in0(and345), .in1(and346), .in2(and347), .in3(and348), .in4(and349), .in5(and350), .in6(and351));
or3$ or_gate24(.out(or24), .in0(and352), .in1(and353), .in2(and354));
or3$ or_gate25(.out(or25), .in0(and355), .in1(and356), .in2(and357));
or5$ or_gate26(.out(or26), .in0(and358), .in1(and359), .in2(and360), .in3(and361), .in4(and362));

assign setd = and0;
assign cleard = and1;
assign size2 = or0;
assign size1 = or1;
assign size0 = or2;
assign op0_2 = or3;
assign op0_1 = or4;
assign op0_0 = or5;
assign op1_2 = or6;
assign op1_1 = or7;
assign op1_0 = or8;
assign op0_reg_4 = and211;
assign op0_reg_3 = or9;
assign op0_reg_2 = or10;
assign op0_reg_1 = or11;
assign op0_reg_0 = or12;
assign op1_reg_4 = and236;
assign op1_reg_3 = or13;
assign op1_reg_2 = or13;
assign op1_reg_1 = or13;
assign op1_reg_0 = or14;
assign alu_op_3 = or15;
assign alu_op_2 = or16;
assign alu_op_1 = or17;
assign alu_op_0 = or18;
assign flag0_2 = or18;
assign flag0_1 = or19;
assign flag0_0 = or20;
assign flag1_2 = or20;
assign flag1_1 = or20;
assign flag1_0 = or21;
assign stack_op_1 = or22;
assign stack_op_0 = or23;
assign rom_control_2 = or24;
assign rom_control_1 = or25;
assign rom_control_0 = or26;
endmodule
