module store_queue();

endmodule
