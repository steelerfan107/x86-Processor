`timescale 1ns / 1ps
module BSF32(in, out, v);
input [31:0] in;
output [31:0] out;
output v; //valid bit

wire in30_not;
wire in29_not;
wire in28_not;
wire in27_not;
wire in26_not;
wire in25_not;
wire in24_not;
wire in23_not;
wire in22_not;
wire in21_not;
wire in20_not;
wire in19_not;
wire in18_not;
wire in17_not;
wire in16_not;
wire in15_not;
wire in14_not;
wire in13_not;
wire in12_not;
wire in11_not;
wire in10_not;
wire in9_not;
wire in8_not;
wire in7_not;
wire in6_not;
wire in5_not;
wire in4_not;
wire in3_not;
wire in2_not;
wire in1_not;
wire in0_not;
wire in30_not_weak;
wire in29_not_weak;
wire in28_not_weak;
wire in27_not_weak;
wire in26_not_weak;
wire in25_not_weak;
wire in24_not_weak;
wire in23_not_weak;
wire in22_not_weak;
wire in21_not_weak;
wire in20_not_weak;
wire in19_not_weak;
wire in18_not_weak;
wire in17_not_weak;
wire in16_not_weak;
wire in15_not_weak;
wire in14_not_weak;
wire in13_not_weak;
wire in12_not_weak;
wire in11_not_weak;
wire in10_not_weak;
wire in9_not_weak;
wire in8_not_weak;
wire in7_not_weak;
wire in6_not_weak;
wire in5_not_weak;
wire in4_not_weak;
wire in3_not_weak;
wire in2_not_weak;
wire in1_not_weak;
wire in0_not_weak;
wire and0;
wire and1;
wire and2;
wire and3;
wire and4;
wire and5;
wire and6;
wire and7;
wire and8;
wire and9;
wire and10;
wire and11;
wire and12;
wire and13;
wire and14;
wire and15;
wire or0;
wire and16;
wire and17;
wire and18;
wire and19;
wire and20;
wire and21;
wire and22;
wire and23;
wire and24;
wire and25;
wire and26;
wire and27;
wire and28;
wire and29;
wire and30;
wire and31;
wire or1;
wire and32;
wire and33;
wire and34;
wire and35;
wire and36;
wire and37;
wire and38;
wire and39;
wire and40;
wire and41;
wire and42;
wire and43;
wire and44;
wire and45;
wire and46;
wire and47;
wire or2;
wire and48;
wire and49;
wire and50;
wire and51;
wire and52;
wire and53;
wire and54;
wire and55;
wire and56;
wire and57;
wire and58;
wire and59;
wire and60;
wire and61;
wire and62;
wire and63;
wire or3;
wire and64;
wire and65;
wire and66;
wire and67;
wire and68;
wire and69;
wire and70;
wire and71;
wire and72;
wire and73;
wire and74;
wire and75;
wire and76;
wire and77;
wire and78;
wire and79;
wire or4;
wire and80;
wire and81;
wire and82;
wire and83;
wire and84;
wire and85;
wire and86;
wire and87;
wire and88;
wire and89;
wire and90;
wire and91;
wire and92;
wire and93;
wire and94;
wire and95;
wire and96;
wire and97;
wire and98;
wire and99;
wire and100;
wire and101;
wire and102;
wire and103;
wire and104;
wire and105;
wire and106;
wire and107;
wire and108;
wire and109;
wire and110;
wire or5;

inv1$ in30_inv (.out(in30_not_weak), .in(in[30]));
inv1$ in29_inv (.out(in29_not_weak), .in(in[29]));
inv1$ in28_inv (.out(in28_not_weak), .in(in[28]));
inv1$ in27_inv (.out(in27_not_weak), .in(in[27]));
inv1$ in26_inv (.out(in26_not_weak), .in(in[26]));
inv1$ in25_inv (.out(in25_not_weak), .in(in[25]));
inv1$ in24_inv (.out(in24_not_weak), .in(in[24]));
inv1$ in23_inv (.out(in23_not_weak), .in(in[23]));
inv1$ in22_inv (.out(in22_not_weak), .in(in[22]));
inv1$ in21_inv (.out(in21_not_weak), .in(in[21]));
inv1$ in20_inv (.out(in20_not_weak), .in(in[20]));
inv1$ in19_inv (.out(in19_not_weak), .in(in[19]));
inv1$ in18_inv (.out(in18_not_weak), .in(in[18]));
inv1$ in17_inv (.out(in17_not_weak), .in(in[17]));
inv1$ in16_inv (.out(in16_not_weak), .in(in[16]));
inv1$ in15_inv (.out(in15_not_weak), .in(in[15]));
inv1$ in14_inv (.out(in14_not_weak), .in(in[14]));
inv1$ in13_inv (.out(in13_not_weak), .in(in[13]));
inv1$ in12_inv (.out(in12_not_weak), .in(in[12]));
inv1$ in11_inv (.out(in11_not_weak), .in(in[11]));
inv1$ in10_inv (.out(in10_not_weak), .in(in[10]));
inv1$ in9_inv (.out(in9_not_weak), .in(in[9]));
inv1$ in8_inv (.out(in8_not_weak), .in(in[8]));
inv1$ in7_inv (.out(in7_not_weak), .in(in[7]));
inv1$ in6_inv (.out(in6_not_weak), .in(in[6]));
inv1$ in5_inv (.out(in5_not_weak), .in(in[5]));
inv1$ in4_inv (.out(in4_not_weak), .in(in[4]));
inv1$ in3_inv (.out(in3_not_weak), .in(in[3]));
inv1$ in2_inv (.out(in2_not_weak), .in(in[2]));
inv1$ in1_inv (.out(in1_not_weak), .in(in[1]));
inv1$ in0_inv (.out(in0_not_weak), .in(in[0]));

bufferH16$ in30_buff(.out(in30_not), .in(in30_not_weak));
bufferH16$ in29_buff(.out(in29_not), .in(in29_not_weak));
bufferH64$ in28_buff(.out(in28_not), .in(in28_not_weak));
bufferH64$ in27_buff(.out(in27_not), .in(in27_not_weak));
bufferH64$ in26_buff(.out(in26_not), .in(in26_not_weak));
bufferH64$ in25_buff(.out(in25_not), .in(in25_not_weak));
bufferH64$ in24_buff(.out(in24_not), .in(in24_not_weak));
bufferH64$ in23_buff(.out(in23_not), .in(in23_not_weak));
bufferH64$ in22_buff(.out(in22_not), .in(in22_not_weak));
bufferH64$ in21_buff(.out(in21_not), .in(in21_not_weak));
bufferH64$ in20_buff(.out(in20_not), .in(in20_not_weak));
bufferH64$ in19_buff(.out(in19_not), .in(in19_not_weak));
bufferH64$ in18_buff(.out(in18_not), .in(in18_not_weak));
bufferH64$ in17_buff(.out(in17_not), .in(in17_not_weak));
bufferH256$ in16_buff(.out(in16_not), .in(in16_not_weak));
bufferH256$ in15_buff(.out(in15_not), .in(in15_not_weak));
bufferH256$ in14_buff(.out(in14_not), .in(in14_not_weak));
bufferH256$ in13_buff(.out(in13_not), .in(in13_not_weak));
bufferH256$ in12_buff(.out(in12_not), .in(in12_not_weak));
bufferH256$ in11_buff(.out(in11_not), .in(in11_not_weak));
bufferH256$ in10_buff(.out(in10_not), .in(in10_not_weak));
bufferH256$ in9_buff(.out(in9_not), .in(in9_not_weak));
bufferH256$ in8_buff(.out(in8_not), .in(in8_not_weak));
bufferH256$ in7_buff(.out(in7_not), .in(in7_not_weak));
bufferH256$ in6_buff(.out(in6_not), .in(in6_not_weak));
bufferH256$ in5_buff(.out(in5_not), .in(in5_not_weak));
bufferH256$ in4_buff(.out(in4_not), .in(in4_not_weak));
bufferH256$ in3_buff(.out(in3_not), .in(in3_not_weak));
bufferH256$ in2_buff(.out(in2_not), .in(in2_not_weak));
bufferH256$ in1_buff(.out(in1_not), .in(in1_not_weak));
bufferH256$ in0_buff(.out(in0_not), .in(in0_not_weak));

and32$ and_gate0(.out(and0), .in0(in[31]), .in1(in30_not), .in2(in29_not), .in3(in28_not), .in4(in27_not), .in5(in26_not), .in6(in25_not), .in7(in24_not), .in8(in23_not), .in9(in22_not), .in10(in21_not), .in11(in20_not), .in12(in19_not), .in13(in18_not), .in14(in17_not), .in15(in16_not), .in16(in15_not), .in17(in14_not), .in18(in13_not), .in19(in12_not), .in20(in11_not), .in21(in10_not), .in22(in9_not), .in23(in8_not), .in24(in7_not), .in25(in6_not), .in26(in5_not), .in27(in4_not), .in28(in3_not), .in29(in2_not), .in30(in1_not), .in31(in0_not));
and31$ and_gate1(.out(and1), .in0(in[30]), .in1(in29_not), .in2(in28_not), .in3(in27_not), .in4(in26_not), .in5(in25_not), .in6(in24_not), .in7(in23_not), .in8(in22_not), .in9(in21_not), .in10(in20_not), .in11(in19_not), .in12(in18_not), .in13(in17_not), .in14(in16_not), .in15(in15_not), .in16(in14_not), .in17(in13_not), .in18(in12_not), .in19(in11_not), .in20(in10_not), .in21(in9_not), .in22(in8_not), .in23(in7_not), .in24(in6_not), .in25(in5_not), .in26(in4_not), .in27(in3_not), .in28(in2_not), .in29(in1_not), .in30(in0_not));
and30$ and_gate2(.out(and2), .in0(in[29]), .in1(in28_not), .in2(in27_not), .in3(in26_not), .in4(in25_not), .in5(in24_not), .in6(in23_not), .in7(in22_not), .in8(in21_not), .in9(in20_not), .in10(in19_not), .in11(in18_not), .in12(in17_not), .in13(in16_not), .in14(in15_not), .in15(in14_not), .in16(in13_not), .in17(in12_not), .in18(in11_not), .in19(in10_not), .in20(in9_not), .in21(in8_not), .in22(in7_not), .in23(in6_not), .in24(in5_not), .in25(in4_not), .in26(in3_not), .in27(in2_not), .in28(in1_not), .in29(in0_not));
and29$ and_gate3(.out(and3), .in0(in[28]), .in1(in27_not), .in2(in26_not), .in3(in25_not), .in4(in24_not), .in5(in23_not), .in6(in22_not), .in7(in21_not), .in8(in20_not), .in9(in19_not), .in10(in18_not), .in11(in17_not), .in12(in16_not), .in13(in15_not), .in14(in14_not), .in15(in13_not), .in16(in12_not), .in17(in11_not), .in18(in10_not), .in19(in9_not), .in20(in8_not), .in21(in7_not), .in22(in6_not), .in23(in5_not), .in24(in4_not), .in25(in3_not), .in26(in2_not), .in27(in1_not), .in28(in0_not));
and28$ and_gate4(.out(and4), .in0(in[27]), .in1(in26_not), .in2(in25_not), .in3(in24_not), .in4(in23_not), .in5(in22_not), .in6(in21_not), .in7(in20_not), .in8(in19_not), .in9(in18_not), .in10(in17_not), .in11(in16_not), .in12(in15_not), .in13(in14_not), .in14(in13_not), .in15(in12_not), .in16(in11_not), .in17(in10_not), .in18(in9_not), .in19(in8_not), .in20(in7_not), .in21(in6_not), .in22(in5_not), .in23(in4_not), .in24(in3_not), .in25(in2_not), .in26(in1_not), .in27(in0_not));
and27$ and_gate5(.out(and5), .in0(in[26]), .in1(in25_not), .in2(in24_not), .in3(in23_not), .in4(in22_not), .in5(in21_not), .in6(in20_not), .in7(in19_not), .in8(in18_not), .in9(in17_not), .in10(in16_not), .in11(in15_not), .in12(in14_not), .in13(in13_not), .in14(in12_not), .in15(in11_not), .in16(in10_not), .in17(in9_not), .in18(in8_not), .in19(in7_not), .in20(in6_not), .in21(in5_not), .in22(in4_not), .in23(in3_not), .in24(in2_not), .in25(in1_not), .in26(in0_not));
and26$ and_gate6(.out(and6), .in0(in[25]), .in1(in24_not), .in2(in23_not), .in3(in22_not), .in4(in21_not), .in5(in20_not), .in6(in19_not), .in7(in18_not), .in8(in17_not), .in9(in16_not), .in10(in15_not), .in11(in14_not), .in12(in13_not), .in13(in12_not), .in14(in11_not), .in15(in10_not), .in16(in9_not), .in17(in8_not), .in18(in7_not), .in19(in6_not), .in20(in5_not), .in21(in4_not), .in22(in3_not), .in23(in2_not), .in24(in1_not), .in25(in0_not));
and25$ and_gate7(.out(and7), .in0(in[24]), .in1(in23_not), .in2(in22_not), .in3(in21_not), .in4(in20_not), .in5(in19_not), .in6(in18_not), .in7(in17_not), .in8(in16_not), .in9(in15_not), .in10(in14_not), .in11(in13_not), .in12(in12_not), .in13(in11_not), .in14(in10_not), .in15(in9_not), .in16(in8_not), .in17(in7_not), .in18(in6_not), .in19(in5_not), .in20(in4_not), .in21(in3_not), .in22(in2_not), .in23(in1_not), .in24(in0_not));
and24$ and_gate8(.out(and8), .in0(in[23]), .in1(in22_not), .in2(in21_not), .in3(in20_not), .in4(in19_not), .in5(in18_not), .in6(in17_not), .in7(in16_not), .in8(in15_not), .in9(in14_not), .in10(in13_not), .in11(in12_not), .in12(in11_not), .in13(in10_not), .in14(in9_not), .in15(in8_not), .in16(in7_not), .in17(in6_not), .in18(in5_not), .in19(in4_not), .in20(in3_not), .in21(in2_not), .in22(in1_not), .in23(in0_not));
and23$ and_gate9(.out(and9), .in0(in[22]), .in1(in21_not), .in2(in20_not), .in3(in19_not), .in4(in18_not), .in5(in17_not), .in6(in16_not), .in7(in15_not), .in8(in14_not), .in9(in13_not), .in10(in12_not), .in11(in11_not), .in12(in10_not), .in13(in9_not), .in14(in8_not), .in15(in7_not), .in16(in6_not), .in17(in5_not), .in18(in4_not), .in19(in3_not), .in20(in2_not), .in21(in1_not), .in22(in0_not));
and22$ and_gate10(.out(and10), .in0(in[21]), .in1(in20_not), .in2(in19_not), .in3(in18_not), .in4(in17_not), .in5(in16_not), .in6(in15_not), .in7(in14_not), .in8(in13_not), .in9(in12_not), .in10(in11_not), .in11(in10_not), .in12(in9_not), .in13(in8_not), .in14(in7_not), .in15(in6_not), .in16(in5_not), .in17(in4_not), .in18(in3_not), .in19(in2_not), .in20(in1_not), .in21(in0_not));
and21$ and_gate11(.out(and11), .in0(in[20]), .in1(in19_not), .in2(in18_not), .in3(in17_not), .in4(in16_not), .in5(in15_not), .in6(in14_not), .in7(in13_not), .in8(in12_not), .in9(in11_not), .in10(in10_not), .in11(in9_not), .in12(in8_not), .in13(in7_not), .in14(in6_not), .in15(in5_not), .in16(in4_not), .in17(in3_not), .in18(in2_not), .in19(in1_not), .in20(in0_not));
and19$ and_gate12(.out(and12), .in0(in[18]), .in1(in17_not), .in2(in16_not), .in3(in15_not), .in4(in14_not), .in5(in13_not), .in6(in12_not), .in7(in11_not), .in8(in10_not), .in9(in9_not), .in10(in8_not), .in11(in7_not), .in12(in6_not), .in13(in5_not), .in14(in4_not), .in15(in3_not), .in16(in2_not), .in17(in1_not), .in18(in0_not));
and20$ and_gate13(.out(and13), .in0(in[19]), .in1(in18_not), .in2(in17_not), .in3(in16_not), .in4(in15_not), .in5(in14_not), .in6(in13_not), .in7(in12_not), .in8(in11_not), .in9(in10_not), .in10(in9_not), .in11(in8_not), .in12(in7_not), .in13(in6_not), .in14(in5_not), .in15(in4_not), .in16(in3_not), .in17(in2_not), .in18(in1_not), .in19(in0_not));
and17$ and_gate14(.out(and14), .in0(in[16]), .in1(in15_not), .in2(in14_not), .in3(in13_not), .in4(in12_not), .in5(in11_not), .in6(in10_not), .in7(in9_not), .in8(in8_not), .in9(in7_not), .in10(in6_not), .in11(in5_not), .in12(in4_not), .in13(in3_not), .in14(in2_not), .in15(in1_not), .in16(in0_not));
and18$ and_gate15(.out(and15), .in0(in[17]), .in1(in16_not), .in2(in15_not), .in3(in14_not), .in4(in13_not), .in5(in12_not), .in6(in11_not), .in7(in10_not), .in8(in9_not), .in9(in8_not), .in10(in7_not), .in11(in6_not), .in12(in5_not), .in13(in4_not), .in14(in3_not), .in15(in2_not), .in16(in1_not), .in17(in0_not));
and32$ and_gate16(.out(and16), .in0(in[31]), .in1(in30_not), .in2(in29_not), .in3(in28_not), .in4(in27_not), .in5(in26_not), .in6(in25_not), .in7(in24_not), .in8(in23_not), .in9(in22_not), .in10(in21_not), .in11(in20_not), .in12(in19_not), .in13(in18_not), .in14(in17_not), .in15(in16_not), .in16(in15_not), .in17(in14_not), .in18(in13_not), .in19(in12_not), .in20(in11_not), .in21(in10_not), .in22(in9_not), .in23(in8_not), .in24(in7_not), .in25(in6_not), .in26(in5_not), .in27(in4_not), .in28(in3_not), .in29(in2_not), .in30(in1_not), .in31(in0_not));
and31$ and_gate17(.out(and17), .in0(in[30]), .in1(in29_not), .in2(in28_not), .in3(in27_not), .in4(in26_not), .in5(in25_not), .in6(in24_not), .in7(in23_not), .in8(in22_not), .in9(in21_not), .in10(in20_not), .in11(in19_not), .in12(in18_not), .in13(in17_not), .in14(in16_not), .in15(in15_not), .in16(in14_not), .in17(in13_not), .in18(in12_not), .in19(in11_not), .in20(in10_not), .in21(in9_not), .in22(in8_not), .in23(in7_not), .in24(in6_not), .in25(in5_not), .in26(in4_not), .in27(in3_not), .in28(in2_not), .in29(in1_not), .in30(in0_not));
and30$ and_gate18(.out(and18), .in0(in[29]), .in1(in28_not), .in2(in27_not), .in3(in26_not), .in4(in25_not), .in5(in24_not), .in6(in23_not), .in7(in22_not), .in8(in21_not), .in9(in20_not), .in10(in19_not), .in11(in18_not), .in12(in17_not), .in13(in16_not), .in14(in15_not), .in15(in14_not), .in16(in13_not), .in17(in12_not), .in18(in11_not), .in19(in10_not), .in20(in9_not), .in21(in8_not), .in22(in7_not), .in23(in6_not), .in24(in5_not), .in25(in4_not), .in26(in3_not), .in27(in2_not), .in28(in1_not), .in29(in0_not));
and29$ and_gate19(.out(and19), .in0(in[28]), .in1(in27_not), .in2(in26_not), .in3(in25_not), .in4(in24_not), .in5(in23_not), .in6(in22_not), .in7(in21_not), .in8(in20_not), .in9(in19_not), .in10(in18_not), .in11(in17_not), .in12(in16_not), .in13(in15_not), .in14(in14_not), .in15(in13_not), .in16(in12_not), .in17(in11_not), .in18(in10_not), .in19(in9_not), .in20(in8_not), .in21(in7_not), .in22(in6_not), .in23(in5_not), .in24(in4_not), .in25(in3_not), .in26(in2_not), .in27(in1_not), .in28(in0_not));
and28$ and_gate20(.out(and20), .in0(in[27]), .in1(in26_not), .in2(in25_not), .in3(in24_not), .in4(in23_not), .in5(in22_not), .in6(in21_not), .in7(in20_not), .in8(in19_not), .in9(in18_not), .in10(in17_not), .in11(in16_not), .in12(in15_not), .in13(in14_not), .in14(in13_not), .in15(in12_not), .in16(in11_not), .in17(in10_not), .in18(in9_not), .in19(in8_not), .in20(in7_not), .in21(in6_not), .in22(in5_not), .in23(in4_not), .in24(in3_not), .in25(in2_not), .in26(in1_not), .in27(in0_not));
and27$ and_gate21(.out(and21), .in0(in[26]), .in1(in25_not), .in2(in24_not), .in3(in23_not), .in4(in22_not), .in5(in21_not), .in6(in20_not), .in7(in19_not), .in8(in18_not), .in9(in17_not), .in10(in16_not), .in11(in15_not), .in12(in14_not), .in13(in13_not), .in14(in12_not), .in15(in11_not), .in16(in10_not), .in17(in9_not), .in18(in8_not), .in19(in7_not), .in20(in6_not), .in21(in5_not), .in22(in4_not), .in23(in3_not), .in24(in2_not), .in25(in1_not), .in26(in0_not));
and26$ and_gate22(.out(and22), .in0(in[25]), .in1(in24_not), .in2(in23_not), .in3(in22_not), .in4(in21_not), .in5(in20_not), .in6(in19_not), .in7(in18_not), .in8(in17_not), .in9(in16_not), .in10(in15_not), .in11(in14_not), .in12(in13_not), .in13(in12_not), .in14(in11_not), .in15(in10_not), .in16(in9_not), .in17(in8_not), .in18(in7_not), .in19(in6_not), .in20(in5_not), .in21(in4_not), .in22(in3_not), .in23(in2_not), .in24(in1_not), .in25(in0_not));
and25$ and_gate23(.out(and23), .in0(in[24]), .in1(in23_not), .in2(in22_not), .in3(in21_not), .in4(in20_not), .in5(in19_not), .in6(in18_not), .in7(in17_not), .in8(in16_not), .in9(in15_not), .in10(in14_not), .in11(in13_not), .in12(in12_not), .in13(in11_not), .in14(in10_not), .in15(in9_not), .in16(in8_not), .in17(in7_not), .in18(in6_not), .in19(in5_not), .in20(in4_not), .in21(in3_not), .in22(in2_not), .in23(in1_not), .in24(in0_not));
and15$ and_gate24(.out(and24), .in0(in[14]), .in1(in13_not), .in2(in12_not), .in3(in11_not), .in4(in10_not), .in5(in9_not), .in6(in8_not), .in7(in7_not), .in8(in6_not), .in9(in5_not), .in10(in4_not), .in11(in3_not), .in12(in2_not), .in13(in1_not), .in14(in0_not));
and13$ and_gate25(.out(and25), .in0(in[12]), .in1(in11_not), .in2(in10_not), .in3(in9_not), .in4(in8_not), .in5(in7_not), .in6(in6_not), .in7(in5_not), .in8(in4_not), .in9(in3_not), .in10(in2_not), .in11(in1_not), .in12(in0_not));
and16$ and_gate26(.out(and26), .in0(in[15]), .in1(in14_not), .in2(in13_not), .in3(in12_not), .in4(in11_not), .in5(in10_not), .in6(in9_not), .in7(in8_not), .in8(in7_not), .in9(in6_not), .in10(in5_not), .in11(in4_not), .in12(in3_not), .in13(in2_not), .in14(in1_not), .in15(in0_not));
and14$ and_gate27(.out(and27), .in0(in[13]), .in1(in12_not), .in2(in11_not), .in3(in10_not), .in4(in9_not), .in5(in8_not), .in6(in7_not), .in7(in6_not), .in8(in5_not), .in9(in4_not), .in10(in3_not), .in11(in2_not), .in12(in1_not), .in13(in0_not));
and11$ and_gate28(.out(and28), .in0(in[10]), .in1(in9_not), .in2(in8_not), .in3(in7_not), .in4(in6_not), .in5(in5_not), .in6(in4_not), .in7(in3_not), .in8(in2_not), .in9(in1_not), .in10(in0_not));
and10$ and_gate29(.out(and29), .in0(in[9]), .in1(in8_not), .in2(in7_not), .in3(in6_not), .in4(in5_not), .in5(in4_not), .in6(in3_not), .in7(in2_not), .in8(in1_not), .in9(in0_not));
and12$ and_gate30(.out(and30), .in0(in[11]), .in1(in10_not), .in2(in9_not), .in3(in8_not), .in4(in7_not), .in5(in6_not), .in6(in5_not), .in7(in4_not), .in8(in3_not), .in9(in2_not), .in10(in1_not), .in11(in0_not));
and9$ and_gate31(.out(and31), .in0(in[8]), .in1(in7_not), .in2(in6_not), .in3(in5_not), .in4(in4_not), .in5(in3_not), .in6(in2_not), .in7(in1_not), .in8(in0_not));
and32$ and_gate32(.out(and32), .in0(in[31]), .in1(in30_not), .in2(in29_not), .in3(in28_not), .in4(in27_not), .in5(in26_not), .in6(in25_not), .in7(in24_not), .in8(in23_not), .in9(in22_not), .in10(in21_not), .in11(in20_not), .in12(in19_not), .in13(in18_not), .in14(in17_not), .in15(in16_not), .in16(in15_not), .in17(in14_not), .in18(in13_not), .in19(in12_not), .in20(in11_not), .in21(in10_not), .in22(in9_not), .in23(in8_not), .in24(in7_not), .in25(in6_not), .in26(in5_not), .in27(in4_not), .in28(in3_not), .in29(in2_not), .in30(in1_not), .in31(in0_not));
and31$ and_gate33(.out(and33), .in0(in[30]), .in1(in29_not), .in2(in28_not), .in3(in27_not), .in4(in26_not), .in5(in25_not), .in6(in24_not), .in7(in23_not), .in8(in22_not), .in9(in21_not), .in10(in20_not), .in11(in19_not), .in12(in18_not), .in13(in17_not), .in14(in16_not), .in15(in15_not), .in16(in14_not), .in17(in13_not), .in18(in12_not), .in19(in11_not), .in20(in10_not), .in21(in9_not), .in22(in8_not), .in23(in7_not), .in24(in6_not), .in25(in5_not), .in26(in4_not), .in27(in3_not), .in28(in2_not), .in29(in1_not), .in30(in0_not));
and30$ and_gate34(.out(and34), .in0(in[29]), .in1(in28_not), .in2(in27_not), .in3(in26_not), .in4(in25_not), .in5(in24_not), .in6(in23_not), .in7(in22_not), .in8(in21_not), .in9(in20_not), .in10(in19_not), .in11(in18_not), .in12(in17_not), .in13(in16_not), .in14(in15_not), .in15(in14_not), .in16(in13_not), .in17(in12_not), .in18(in11_not), .in19(in10_not), .in20(in9_not), .in21(in8_not), .in22(in7_not), .in23(in6_not), .in24(in5_not), .in25(in4_not), .in26(in3_not), .in27(in2_not), .in28(in1_not), .in29(in0_not));
and29$ and_gate35(.out(and35), .in0(in[28]), .in1(in27_not), .in2(in26_not), .in3(in25_not), .in4(in24_not), .in5(in23_not), .in6(in22_not), .in7(in21_not), .in8(in20_not), .in9(in19_not), .in10(in18_not), .in11(in17_not), .in12(in16_not), .in13(in15_not), .in14(in14_not), .in15(in13_not), .in16(in12_not), .in17(in11_not), .in18(in10_not), .in19(in9_not), .in20(in8_not), .in21(in7_not), .in22(in6_not), .in23(in5_not), .in24(in4_not), .in25(in3_not), .in26(in2_not), .in27(in1_not), .in28(in0_not));
and24$ and_gate36(.out(and36), .in0(in[23]), .in1(in22_not), .in2(in21_not), .in3(in20_not), .in4(in19_not), .in5(in18_not), .in6(in17_not), .in7(in16_not), .in8(in15_not), .in9(in14_not), .in10(in13_not), .in11(in12_not), .in12(in11_not), .in13(in10_not), .in14(in9_not), .in15(in8_not), .in16(in7_not), .in17(in6_not), .in18(in5_not), .in19(in4_not), .in20(in3_not), .in21(in2_not), .in22(in1_not), .in23(in0_not));
and23$ and_gate37(.out(and37), .in0(in[22]), .in1(in21_not), .in2(in20_not), .in3(in19_not), .in4(in18_not), .in5(in17_not), .in6(in16_not), .in7(in15_not), .in8(in14_not), .in9(in13_not), .in10(in12_not), .in11(in11_not), .in12(in10_not), .in13(in9_not), .in14(in8_not), .in15(in7_not), .in16(in6_not), .in17(in5_not), .in18(in4_not), .in19(in3_not), .in20(in2_not), .in21(in1_not), .in22(in0_not));
and22$ and_gate38(.out(and38), .in0(in[21]), .in1(in20_not), .in2(in19_not), .in3(in18_not), .in4(in17_not), .in5(in16_not), .in6(in15_not), .in7(in14_not), .in8(in13_not), .in9(in12_not), .in10(in11_not), .in11(in10_not), .in12(in9_not), .in13(in8_not), .in14(in7_not), .in15(in6_not), .in16(in5_not), .in17(in4_not), .in18(in3_not), .in19(in2_not), .in20(in1_not), .in21(in0_not));
and21$ and_gate39(.out(and39), .in0(in[20]), .in1(in19_not), .in2(in18_not), .in3(in17_not), .in4(in16_not), .in5(in15_not), .in6(in14_not), .in7(in13_not), .in8(in12_not), .in9(in11_not), .in10(in10_not), .in11(in9_not), .in12(in8_not), .in13(in7_not), .in14(in6_not), .in15(in5_not), .in16(in4_not), .in17(in3_not), .in18(in2_not), .in19(in1_not), .in20(in0_not));
and15$ and_gate40(.out(and40), .in0(in[14]), .in1(in13_not), .in2(in12_not), .in3(in11_not), .in4(in10_not), .in5(in9_not), .in6(in8_not), .in7(in7_not), .in8(in6_not), .in9(in5_not), .in10(in4_not), .in11(in3_not), .in12(in2_not), .in13(in1_not), .in14(in0_not));
and13$ and_gate41(.out(and41), .in0(in[12]), .in1(in11_not), .in2(in10_not), .in3(in9_not), .in4(in8_not), .in5(in7_not), .in6(in6_not), .in7(in5_not), .in8(in4_not), .in9(in3_not), .in10(in2_not), .in11(in1_not), .in12(in0_not));
and16$ and_gate42(.out(and42), .in0(in[15]), .in1(in14_not), .in2(in13_not), .in3(in12_not), .in4(in11_not), .in5(in10_not), .in6(in9_not), .in7(in8_not), .in8(in7_not), .in9(in6_not), .in10(in5_not), .in11(in4_not), .in12(in3_not), .in13(in2_not), .in14(in1_not), .in15(in0_not));
and14$ and_gate43(.out(and43), .in0(in[13]), .in1(in12_not), .in2(in11_not), .in3(in10_not), .in4(in9_not), .in5(in8_not), .in6(in7_not), .in7(in6_not), .in8(in5_not), .in9(in4_not), .in10(in3_not), .in11(in2_not), .in12(in1_not), .in13(in0_not));
and7$ and_gate44(.out(and44), .in0(in[6]), .in1(in5_not), .in2(in4_not), .in3(in3_not), .in4(in2_not), .in5(in1_not), .in6(in0_not));
and6$ and_gate45(.out(and45), .in0(in[5]), .in1(in4_not), .in2(in3_not), .in3(in2_not), .in4(in1_not), .in5(in0_not));
and8$ and_gate46(.out(and46), .in0(in[7]), .in1(in6_not), .in2(in5_not), .in3(in4_not), .in4(in3_not), .in5(in2_not), .in6(in1_not), .in7(in0_not));
and5$ and_gate47(.out(and47), .in0(in[4]), .in1(in3_not), .in2(in2_not), .in3(in1_not), .in4(in0_not));
and32$ and_gate48(.out(and48), .in0(in[31]), .in1(in30_not), .in2(in29_not), .in3(in28_not), .in4(in27_not), .in5(in26_not), .in6(in25_not), .in7(in24_not), .in8(in23_not), .in9(in22_not), .in10(in21_not), .in11(in20_not), .in12(in19_not), .in13(in18_not), .in14(in17_not), .in15(in16_not), .in16(in15_not), .in17(in14_not), .in18(in13_not), .in19(in12_not), .in20(in11_not), .in21(in10_not), .in22(in9_not), .in23(in8_not), .in24(in7_not), .in25(in6_not), .in26(in5_not), .in27(in4_not), .in28(in3_not), .in29(in2_not), .in30(in1_not), .in31(in0_not));
and31$ and_gate49(.out(and49), .in0(in[30]), .in1(in29_not), .in2(in28_not), .in3(in27_not), .in4(in26_not), .in5(in25_not), .in6(in24_not), .in7(in23_not), .in8(in22_not), .in9(in21_not), .in10(in20_not), .in11(in19_not), .in12(in18_not), .in13(in17_not), .in14(in16_not), .in15(in15_not), .in16(in14_not), .in17(in13_not), .in18(in12_not), .in19(in11_not), .in20(in10_not), .in21(in9_not), .in22(in8_not), .in23(in7_not), .in24(in6_not), .in25(in5_not), .in26(in4_not), .in27(in3_not), .in28(in2_not), .in29(in1_not), .in30(in0_not));
and28$ and_gate50(.out(and50), .in0(in[27]), .in1(in26_not), .in2(in25_not), .in3(in24_not), .in4(in23_not), .in5(in22_not), .in6(in21_not), .in7(in20_not), .in8(in19_not), .in9(in18_not), .in10(in17_not), .in11(in16_not), .in12(in15_not), .in13(in14_not), .in14(in13_not), .in15(in12_not), .in16(in11_not), .in17(in10_not), .in18(in9_not), .in19(in8_not), .in20(in7_not), .in21(in6_not), .in22(in5_not), .in23(in4_not), .in24(in3_not), .in25(in2_not), .in26(in1_not), .in27(in0_not));
and27$ and_gate51(.out(and51), .in0(in[26]), .in1(in25_not), .in2(in24_not), .in3(in23_not), .in4(in22_not), .in5(in21_not), .in6(in20_not), .in7(in19_not), .in8(in18_not), .in9(in17_not), .in10(in16_not), .in11(in15_not), .in12(in14_not), .in13(in13_not), .in14(in12_not), .in15(in11_not), .in16(in10_not), .in17(in9_not), .in18(in8_not), .in19(in7_not), .in20(in6_not), .in21(in5_not), .in22(in4_not), .in23(in3_not), .in24(in2_not), .in25(in1_not), .in26(in0_not));
and24$ and_gate52(.out(and52), .in0(in[23]), .in1(in22_not), .in2(in21_not), .in3(in20_not), .in4(in19_not), .in5(in18_not), .in6(in17_not), .in7(in16_not), .in8(in15_not), .in9(in14_not), .in10(in13_not), .in11(in12_not), .in12(in11_not), .in13(in10_not), .in14(in9_not), .in15(in8_not), .in16(in7_not), .in17(in6_not), .in18(in5_not), .in19(in4_not), .in20(in3_not), .in21(in2_not), .in22(in1_not), .in23(in0_not));
and23$ and_gate53(.out(and53), .in0(in[22]), .in1(in21_not), .in2(in20_not), .in3(in19_not), .in4(in18_not), .in5(in17_not), .in6(in16_not), .in7(in15_not), .in8(in14_not), .in9(in13_not), .in10(in12_not), .in11(in11_not), .in12(in10_not), .in13(in9_not), .in14(in8_not), .in15(in7_not), .in16(in6_not), .in17(in5_not), .in18(in4_not), .in19(in3_not), .in20(in2_not), .in21(in1_not), .in22(in0_not));
and19$ and_gate54(.out(and54), .in0(in[18]), .in1(in17_not), .in2(in16_not), .in3(in15_not), .in4(in14_not), .in5(in13_not), .in6(in12_not), .in7(in11_not), .in8(in10_not), .in9(in9_not), .in10(in8_not), .in11(in7_not), .in12(in6_not), .in13(in5_not), .in14(in4_not), .in15(in3_not), .in16(in2_not), .in17(in1_not), .in18(in0_not));
and20$ and_gate55(.out(and55), .in0(in[19]), .in1(in18_not), .in2(in17_not), .in3(in16_not), .in4(in15_not), .in5(in14_not), .in6(in13_not), .in7(in12_not), .in8(in11_not), .in9(in10_not), .in10(in9_not), .in11(in8_not), .in12(in7_not), .in13(in6_not), .in14(in5_not), .in15(in4_not), .in16(in3_not), .in17(in2_not), .in18(in1_not), .in19(in0_not));
and15$ and_gate56(.out(and56), .in0(in[14]), .in1(in13_not), .in2(in12_not), .in3(in11_not), .in4(in10_not), .in5(in9_not), .in6(in8_not), .in7(in7_not), .in8(in6_not), .in9(in5_not), .in10(in4_not), .in11(in3_not), .in12(in2_not), .in13(in1_not), .in14(in0_not));
and16$ and_gate57(.out(and57), .in0(in[15]), .in1(in14_not), .in2(in13_not), .in3(in12_not), .in4(in11_not), .in5(in10_not), .in6(in9_not), .in7(in8_not), .in8(in7_not), .in9(in6_not), .in10(in5_not), .in11(in4_not), .in12(in3_not), .in13(in2_not), .in14(in1_not), .in15(in0_not));
and11$ and_gate58(.out(and58), .in0(in[10]), .in1(in9_not), .in2(in8_not), .in3(in7_not), .in4(in6_not), .in5(in5_not), .in6(in4_not), .in7(in3_not), .in8(in2_not), .in9(in1_not), .in10(in0_not));
and12$ and_gate59(.out(and59), .in0(in[11]), .in1(in10_not), .in2(in9_not), .in3(in8_not), .in4(in7_not), .in5(in6_not), .in6(in5_not), .in7(in4_not), .in8(in3_not), .in9(in2_not), .in10(in1_not), .in11(in0_not));
and7$ and_gate60(.out(and60), .in0(in[6]), .in1(in5_not), .in2(in4_not), .in3(in3_not), .in4(in2_not), .in5(in1_not), .in6(in0_not));
and4$ and_gate61(.out(and61), .in0(in[3]), .in1(in2_not), .in2(in1_not), .in3(in0_not));
and8$ and_gate62(.out(and62), .in0(in[7]), .in1(in6_not), .in2(in5_not), .in3(in4_not), .in4(in3_not), .in5(in2_not), .in6(in1_not), .in7(in0_not));
and3$ and_gate63(.out(and63), .in0(in[2]), .in1(in1_not), .in2(in0_not));
and32$ and_gate64(.out(and64), .in0(in[31]), .in1(in30_not), .in2(in29_not), .in3(in28_not), .in4(in27_not), .in5(in26_not), .in6(in25_not), .in7(in24_not), .in8(in23_not), .in9(in22_not), .in10(in21_not), .in11(in20_not), .in12(in19_not), .in13(in18_not), .in14(in17_not), .in15(in16_not), .in16(in15_not), .in17(in14_not), .in18(in13_not), .in19(in12_not), .in20(in11_not), .in21(in10_not), .in22(in9_not), .in23(in8_not), .in24(in7_not), .in25(in6_not), .in26(in5_not), .in27(in4_not), .in28(in3_not), .in29(in2_not), .in30(in1_not), .in31(in0_not));
and30$ and_gate65(.out(and65), .in0(in[29]), .in1(in28_not), .in2(in27_not), .in3(in26_not), .in4(in25_not), .in5(in24_not), .in6(in23_not), .in7(in22_not), .in8(in21_not), .in9(in20_not), .in10(in19_not), .in11(in18_not), .in12(in17_not), .in13(in16_not), .in14(in15_not), .in15(in14_not), .in16(in13_not), .in17(in12_not), .in18(in11_not), .in19(in10_not), .in20(in9_not), .in21(in8_not), .in22(in7_not), .in23(in6_not), .in24(in5_not), .in25(in4_not), .in26(in3_not), .in27(in2_not), .in28(in1_not), .in29(in0_not));
and28$ and_gate66(.out(and66), .in0(in[27]), .in1(in26_not), .in2(in25_not), .in3(in24_not), .in4(in23_not), .in5(in22_not), .in6(in21_not), .in7(in20_not), .in8(in19_not), .in9(in18_not), .in10(in17_not), .in11(in16_not), .in12(in15_not), .in13(in14_not), .in14(in13_not), .in15(in12_not), .in16(in11_not), .in17(in10_not), .in18(in9_not), .in19(in8_not), .in20(in7_not), .in21(in6_not), .in22(in5_not), .in23(in4_not), .in24(in3_not), .in25(in2_not), .in26(in1_not), .in27(in0_not));
and26$ and_gate67(.out(and67), .in0(in[25]), .in1(in24_not), .in2(in23_not), .in3(in22_not), .in4(in21_not), .in5(in20_not), .in6(in19_not), .in7(in18_not), .in8(in17_not), .in9(in16_not), .in10(in15_not), .in11(in14_not), .in12(in13_not), .in13(in12_not), .in14(in11_not), .in15(in10_not), .in16(in9_not), .in17(in8_not), .in18(in7_not), .in19(in6_not), .in20(in5_not), .in21(in4_not), .in22(in3_not), .in23(in2_not), .in24(in1_not), .in25(in0_not));
and24$ and_gate68(.out(and68), .in0(in[23]), .in1(in22_not), .in2(in21_not), .in3(in20_not), .in4(in19_not), .in5(in18_not), .in6(in17_not), .in7(in16_not), .in8(in15_not), .in9(in14_not), .in10(in13_not), .in11(in12_not), .in12(in11_not), .in13(in10_not), .in14(in9_not), .in15(in8_not), .in16(in7_not), .in17(in6_not), .in18(in5_not), .in19(in4_not), .in20(in3_not), .in21(in2_not), .in22(in1_not), .in23(in0_not));
and22$ and_gate69(.out(and69), .in0(in[21]), .in1(in20_not), .in2(in19_not), .in3(in18_not), .in4(in17_not), .in5(in16_not), .in6(in15_not), .in7(in14_not), .in8(in13_not), .in9(in12_not), .in10(in11_not), .in11(in10_not), .in12(in9_not), .in13(in8_not), .in14(in7_not), .in15(in6_not), .in16(in5_not), .in17(in4_not), .in18(in3_not), .in19(in2_not), .in20(in1_not), .in21(in0_not));
and20$ and_gate70(.out(and70), .in0(in[19]), .in1(in18_not), .in2(in17_not), .in3(in16_not), .in4(in15_not), .in5(in14_not), .in6(in13_not), .in7(in12_not), .in8(in11_not), .in9(in10_not), .in10(in9_not), .in11(in8_not), .in12(in7_not), .in13(in6_not), .in14(in5_not), .in15(in4_not), .in16(in3_not), .in17(in2_not), .in18(in1_not), .in19(in0_not));
and18$ and_gate71(.out(and71), .in0(in[17]), .in1(in16_not), .in2(in15_not), .in3(in14_not), .in4(in13_not), .in5(in12_not), .in6(in11_not), .in7(in10_not), .in8(in9_not), .in9(in8_not), .in10(in7_not), .in11(in6_not), .in12(in5_not), .in13(in4_not), .in14(in3_not), .in15(in2_not), .in16(in1_not), .in17(in0_not));
and16$ and_gate72(.out(and72), .in0(in[15]), .in1(in14_not), .in2(in13_not), .in3(in12_not), .in4(in11_not), .in5(in10_not), .in6(in9_not), .in7(in8_not), .in8(in7_not), .in9(in6_not), .in10(in5_not), .in11(in4_not), .in12(in3_not), .in13(in2_not), .in14(in1_not), .in15(in0_not));
and14$ and_gate73(.out(and73), .in0(in[13]), .in1(in12_not), .in2(in11_not), .in3(in10_not), .in4(in9_not), .in5(in8_not), .in6(in7_not), .in7(in6_not), .in8(in5_not), .in9(in4_not), .in10(in3_not), .in11(in2_not), .in12(in1_not), .in13(in0_not));
and10$ and_gate74(.out(and74), .in0(in[9]), .in1(in8_not), .in2(in7_not), .in3(in6_not), .in4(in5_not), .in5(in4_not), .in6(in3_not), .in7(in2_not), .in8(in1_not), .in9(in0_not));
and12$ and_gate75(.out(and75), .in0(in[11]), .in1(in10_not), .in2(in9_not), .in3(in8_not), .in4(in7_not), .in5(in6_not), .in6(in5_not), .in7(in4_not), .in8(in3_not), .in9(in2_not), .in10(in1_not), .in11(in0_not));
and6$ and_gate76(.out(and76), .in0(in[5]), .in1(in4_not), .in2(in3_not), .in3(in2_not), .in4(in1_not), .in5(in0_not));
and4$ and_gate77(.out(and77), .in0(in[3]), .in1(in2_not), .in2(in1_not), .in3(in0_not));
and8$ and_gate78(.out(and78), .in0(in[7]), .in1(in6_not), .in2(in5_not), .in3(in4_not), .in4(in3_not), .in5(in2_not), .in6(in1_not), .in7(in0_not));
and2$ and_gate79(.out(and79), .in0(in[1]), .in1(in0_not));
and32$ and_gate80(.out(and80), .in0(in[31]), .in1(in30_not), .in2(in29_not), .in3(in28_not), .in4(in27_not), .in5(in26_not), .in6(in25_not), .in7(in24_not), .in8(in23_not), .in9(in22_not), .in10(in21_not), .in11(in20_not), .in12(in19_not), .in13(in18_not), .in14(in17_not), .in15(in16_not), .in16(in15_not), .in17(in14_not), .in18(in13_not), .in19(in12_not), .in20(in11_not), .in21(in10_not), .in22(in9_not), .in23(in8_not), .in24(in7_not), .in25(in6_not), .in26(in5_not), .in27(in4_not), .in28(in3_not), .in29(in2_not), .in30(in1_not), .in31(in0_not));
and31$ and_gate81(.out(and81), .in0(in[30]), .in1(in29_not), .in2(in28_not), .in3(in27_not), .in4(in26_not), .in5(in25_not), .in6(in24_not), .in7(in23_not), .in8(in22_not), .in9(in21_not), .in10(in20_not), .in11(in19_not), .in12(in18_not), .in13(in17_not), .in14(in16_not), .in15(in15_not), .in16(in14_not), .in17(in13_not), .in18(in12_not), .in19(in11_not), .in20(in10_not), .in21(in9_not), .in22(in8_not), .in23(in7_not), .in24(in6_not), .in25(in5_not), .in26(in4_not), .in27(in3_not), .in28(in2_not), .in29(in1_not), .in30(in0_not));
and30$ and_gate82(.out(and82), .in0(in[29]), .in1(in28_not), .in2(in27_not), .in3(in26_not), .in4(in25_not), .in5(in24_not), .in6(in23_not), .in7(in22_not), .in8(in21_not), .in9(in20_not), .in10(in19_not), .in11(in18_not), .in12(in17_not), .in13(in16_not), .in14(in15_not), .in15(in14_not), .in16(in13_not), .in17(in12_not), .in18(in11_not), .in19(in10_not), .in20(in9_not), .in21(in8_not), .in22(in7_not), .in23(in6_not), .in24(in5_not), .in25(in4_not), .in26(in3_not), .in27(in2_not), .in28(in1_not), .in29(in0_not));
and29$ and_gate83(.out(and83), .in0(in[28]), .in1(in27_not), .in2(in26_not), .in3(in25_not), .in4(in24_not), .in5(in23_not), .in6(in22_not), .in7(in21_not), .in8(in20_not), .in9(in19_not), .in10(in18_not), .in11(in17_not), .in12(in16_not), .in13(in15_not), .in14(in14_not), .in15(in13_not), .in16(in12_not), .in17(in11_not), .in18(in10_not), .in19(in9_not), .in20(in8_not), .in21(in7_not), .in22(in6_not), .in23(in5_not), .in24(in4_not), .in25(in3_not), .in26(in2_not), .in27(in1_not), .in28(in0_not));
and28$ and_gate84(.out(and84), .in0(in[27]), .in1(in26_not), .in2(in25_not), .in3(in24_not), .in4(in23_not), .in5(in22_not), .in6(in21_not), .in7(in20_not), .in8(in19_not), .in9(in18_not), .in10(in17_not), .in11(in16_not), .in12(in15_not), .in13(in14_not), .in14(in13_not), .in15(in12_not), .in16(in11_not), .in17(in10_not), .in18(in9_not), .in19(in8_not), .in20(in7_not), .in21(in6_not), .in22(in5_not), .in23(in4_not), .in24(in3_not), .in25(in2_not), .in26(in1_not), .in27(in0_not));
and27$ and_gate85(.out(and85), .in0(in[26]), .in1(in25_not), .in2(in24_not), .in3(in23_not), .in4(in22_not), .in5(in21_not), .in6(in20_not), .in7(in19_not), .in8(in18_not), .in9(in17_not), .in10(in16_not), .in11(in15_not), .in12(in14_not), .in13(in13_not), .in14(in12_not), .in15(in11_not), .in16(in10_not), .in17(in9_not), .in18(in8_not), .in19(in7_not), .in20(in6_not), .in21(in5_not), .in22(in4_not), .in23(in3_not), .in24(in2_not), .in25(in1_not), .in26(in0_not));
and26$ and_gate86(.out(and86), .in0(in[25]), .in1(in24_not), .in2(in23_not), .in3(in22_not), .in4(in21_not), .in5(in20_not), .in6(in19_not), .in7(in18_not), .in8(in17_not), .in9(in16_not), .in10(in15_not), .in11(in14_not), .in12(in13_not), .in13(in12_not), .in14(in11_not), .in15(in10_not), .in16(in9_not), .in17(in8_not), .in18(in7_not), .in19(in6_not), .in20(in5_not), .in21(in4_not), .in22(in3_not), .in23(in2_not), .in24(in1_not), .in25(in0_not));
and25$ and_gate87(.out(and87), .in0(in[24]), .in1(in23_not), .in2(in22_not), .in3(in21_not), .in4(in20_not), .in5(in19_not), .in6(in18_not), .in7(in17_not), .in8(in16_not), .in9(in15_not), .in10(in14_not), .in11(in13_not), .in12(in12_not), .in13(in11_not), .in14(in10_not), .in15(in9_not), .in16(in8_not), .in17(in7_not), .in18(in6_not), .in19(in5_not), .in20(in4_not), .in21(in3_not), .in22(in2_not), .in23(in1_not), .in24(in0_not));
and24$ and_gate88(.out(and88), .in0(in[23]), .in1(in22_not), .in2(in21_not), .in3(in20_not), .in4(in19_not), .in5(in18_not), .in6(in17_not), .in7(in16_not), .in8(in15_not), .in9(in14_not), .in10(in13_not), .in11(in12_not), .in12(in11_not), .in13(in10_not), .in14(in9_not), .in15(in8_not), .in16(in7_not), .in17(in6_not), .in18(in5_not), .in19(in4_not), .in20(in3_not), .in21(in2_not), .in22(in1_not), .in23(in0_not));
and23$ and_gate89(.out(and89), .in0(in[22]), .in1(in21_not), .in2(in20_not), .in3(in19_not), .in4(in18_not), .in5(in17_not), .in6(in16_not), .in7(in15_not), .in8(in14_not), .in9(in13_not), .in10(in12_not), .in11(in11_not), .in12(in10_not), .in13(in9_not), .in14(in8_not), .in15(in7_not), .in16(in6_not), .in17(in5_not), .in18(in4_not), .in19(in3_not), .in20(in2_not), .in21(in1_not), .in22(in0_not));
and22$ and_gate90(.out(and90), .in0(in[21]), .in1(in20_not), .in2(in19_not), .in3(in18_not), .in4(in17_not), .in5(in16_not), .in6(in15_not), .in7(in14_not), .in8(in13_not), .in9(in12_not), .in10(in11_not), .in11(in10_not), .in12(in9_not), .in13(in8_not), .in14(in7_not), .in15(in6_not), .in16(in5_not), .in17(in4_not), .in18(in3_not), .in19(in2_not), .in20(in1_not), .in21(in0_not));
and21$ and_gate91(.out(and91), .in0(in[20]), .in1(in19_not), .in2(in18_not), .in3(in17_not), .in4(in16_not), .in5(in15_not), .in6(in14_not), .in7(in13_not), .in8(in12_not), .in9(in11_not), .in10(in10_not), .in11(in9_not), .in12(in8_not), .in13(in7_not), .in14(in6_not), .in15(in5_not), .in16(in4_not), .in17(in3_not), .in18(in2_not), .in19(in1_not), .in20(in0_not));
and19$ and_gate92(.out(and92), .in0(in[18]), .in1(in17_not), .in2(in16_not), .in3(in15_not), .in4(in14_not), .in5(in13_not), .in6(in12_not), .in7(in11_not), .in8(in10_not), .in9(in9_not), .in10(in8_not), .in11(in7_not), .in12(in6_not), .in13(in5_not), .in14(in4_not), .in15(in3_not), .in16(in2_not), .in17(in1_not), .in18(in0_not));
and20$ and_gate93(.out(and93), .in0(in[19]), .in1(in18_not), .in2(in17_not), .in3(in16_not), .in4(in15_not), .in5(in14_not), .in6(in13_not), .in7(in12_not), .in8(in11_not), .in9(in10_not), .in10(in9_not), .in11(in8_not), .in12(in7_not), .in13(in6_not), .in14(in5_not), .in15(in4_not), .in16(in3_not), .in17(in2_not), .in18(in1_not), .in19(in0_not));
and17$ and_gate94(.out(and94), .in0(in[16]), .in1(in15_not), .in2(in14_not), .in3(in13_not), .in4(in12_not), .in5(in11_not), .in6(in10_not), .in7(in9_not), .in8(in8_not), .in9(in7_not), .in10(in6_not), .in11(in5_not), .in12(in4_not), .in13(in3_not), .in14(in2_not), .in15(in1_not), .in16(in0_not));
and18$ and_gate95(.out(and95), .in0(in[17]), .in1(in16_not), .in2(in15_not), .in3(in14_not), .in4(in13_not), .in5(in12_not), .in6(in11_not), .in7(in10_not), .in8(in9_not), .in9(in8_not), .in10(in7_not), .in11(in6_not), .in12(in5_not), .in13(in4_not), .in14(in3_not), .in15(in2_not), .in16(in1_not), .in17(in0_not));
and15$ and_gate96(.out(and96), .in0(in[14]), .in1(in13_not), .in2(in12_not), .in3(in11_not), .in4(in10_not), .in5(in9_not), .in6(in8_not), .in7(in7_not), .in8(in6_not), .in9(in5_not), .in10(in4_not), .in11(in3_not), .in12(in2_not), .in13(in1_not), .in14(in0_not));
and13$ and_gate97(.out(and97), .in0(in[12]), .in1(in11_not), .in2(in10_not), .in3(in9_not), .in4(in8_not), .in5(in7_not), .in6(in6_not), .in7(in5_not), .in8(in4_not), .in9(in3_not), .in10(in2_not), .in11(in1_not), .in12(in0_not));
and16$ and_gate98(.out(and98), .in0(in[15]), .in1(in14_not), .in2(in13_not), .in3(in12_not), .in4(in11_not), .in5(in10_not), .in6(in9_not), .in7(in8_not), .in8(in7_not), .in9(in6_not), .in10(in5_not), .in11(in4_not), .in12(in3_not), .in13(in2_not), .in14(in1_not), .in15(in0_not));
and14$ and_gate99(.out(and99), .in0(in[13]), .in1(in12_not), .in2(in11_not), .in3(in10_not), .in4(in9_not), .in5(in8_not), .in6(in7_not), .in7(in6_not), .in8(in5_not), .in9(in4_not), .in10(in3_not), .in11(in2_not), .in12(in1_not), .in13(in0_not));
and11$ and_gate100(.out(and100), .in0(in[10]), .in1(in9_not), .in2(in8_not), .in3(in7_not), .in4(in6_not), .in5(in5_not), .in6(in4_not), .in7(in3_not), .in8(in2_not), .in9(in1_not), .in10(in0_not));
and10$ and_gate101(.out(and101), .in0(in[9]), .in1(in8_not), .in2(in7_not), .in3(in6_not), .in4(in5_not), .in5(in4_not), .in6(in3_not), .in7(in2_not), .in8(in1_not), .in9(in0_not));
and12$ and_gate102(.out(and102), .in0(in[11]), .in1(in10_not), .in2(in9_not), .in3(in8_not), .in4(in7_not), .in5(in6_not), .in6(in5_not), .in7(in4_not), .in8(in3_not), .in9(in2_not), .in10(in1_not), .in11(in0_not));
and7$ and_gate103(.out(and103), .in0(in[6]), .in1(in5_not), .in2(in4_not), .in3(in3_not), .in4(in2_not), .in5(in1_not), .in6(in0_not));
and6$ and_gate104(.out(and104), .in0(in[5]), .in1(in4_not), .in2(in3_not), .in3(in2_not), .in4(in1_not), .in5(in0_not));
and4$ and_gate105(.out(and105), .in0(in[3]), .in1(in2_not), .in2(in1_not), .in3(in0_not));
and8$ and_gate106(.out(and106), .in0(in[7]), .in1(in6_not), .in2(in5_not), .in3(in4_not), .in4(in3_not), .in5(in2_not), .in6(in1_not), .in7(in0_not));
and9$ and_gate107(.out(and107), .in0(in[8]), .in1(in7_not), .in2(in6_not), .in3(in5_not), .in4(in4_not), .in5(in3_not), .in6(in2_not), .in7(in1_not), .in8(in0_not));
and5$ and_gate108(.out(and108), .in0(in[4]), .in1(in3_not), .in2(in2_not), .in3(in1_not), .in4(in0_not));
and3$ and_gate109(.out(and109), .in0(in[2]), .in1(in1_not), .in2(in0_not));
and2$ and_gate110(.out(and110), .in0(in[1]), .in1(in0_not));

or16$ or_gate0(.out(or0), .in0(and0), .in1(and1), .in2(and2), .in3(and3), .in4(and4), .in5(and5), .in6(and6), .in7(and7), .in8(and8), .in9(and9), .in10(and10), .in11(and11), .in12(and12), .in13(and13), .in14(and14), .in15(and15));
or16$ or_gate1(.out(or1), .in0(and16), .in1(and17), .in2(and18), .in3(and19), .in4(and20), .in5(and21), .in6(and22), .in7(and23), .in8(and24), .in9(and25), .in10(and26), .in11(and27), .in12(and28), .in13(and29), .in14(and30), .in15(and31));
or16$ or_gate2(.out(or2), .in0(and32), .in1(and33), .in2(and34), .in3(and35), .in4(and36), .in5(and37), .in6(and38), .in7(and39), .in8(and40), .in9(and41), .in10(and42), .in11(and43), .in12(and44), .in13(and45), .in14(and46), .in15(and47));
or16$ or_gate3(.out(or3), .in0(and48), .in1(and49), .in2(and50), .in3(and51), .in4(and52), .in5(and53), .in6(and54), .in7(and55), .in8(and56), .in9(and57), .in10(and58), .in11(and59), .in12(and60), .in13(and61), .in14(and62), .in15(and63));
or16$ or_gate4(.out(or4), .in0(and64), .in1(and65), .in2(and66), .in3(and67), .in4(and68), .in5(and69), .in6(and70), .in7(and71), .in8(and72), .in9(and73), .in10(and74), .in11(and75), .in12(and76), .in13(and77), .in14(and78), .in15(and79));
or32$ or_gate5(.out(or5), .in0(and80), .in1(and81), .in2(and82), .in3(and83), .in4(and84), .in5(and85), .in6(and86), .in7(and87), .in8(and88), .in9(and89), .in10(and90), .in11(and91), .in12(and92), .in13(and93), .in14(and94), .in15(and95), .in16(and96), .in17(and97), .in18(and98), .in19(and99), .in20(and100), .in21(and101), .in22(and102), .in23(and103), .in24(and104), .in25(and105), .in26(and106), .in27(and107), .in28(in[0]), .in29(and108), .in30(and109), .in31(and110));

assign out[4] = or0;
assign out[3] = or1;
assign out[2] = or2;
assign out[1] = or3;
assign out[0] = or4;
assign v = or5;

assign out[31:5] = 27'h0000000;

endmodule

`timescale 1ns / 1ps
module BSF16(in, out, v);
input [15:0] in;
output [31:0] out;
output v;

wire in14_not;
wire in13_not;
wire in12_not;
wire in11_not;
wire in10_not;
wire in9_not;
wire in8_not;
wire in7_not;
wire in6_not;
wire in5_not;
wire in4_not;
wire in3_not;
wire in2_not;
wire in1_not;
wire in0_not;
wire in14_not_weak;
wire in13_not_weak;
wire in12_not_weak;
wire in11_not_weak;
wire in10_not_weak;
wire in9_not_weak;
wire in8_not_weak;
wire in7_not_weak;
wire in6_not_weak;
wire in5_not_weak;
wire in4_not_weak;
wire in3_not_weak;
wire in2_not_weak;
wire in1_not_weak;
wire in0_not_weak;
wire and0;
wire and1;
wire and2;
wire and3;
wire and4;
wire and5;
wire and6;
wire and7;
wire or0;
wire and8;
wire and9;
wire and10;
wire and11;
wire and12;
wire and13;
wire and14;
wire and15;
wire or1;
wire and16;
wire and17;
wire and18;
wire and19;
wire and20;
wire and21;
wire and22;
wire and23;
wire or2;
wire and24;
wire and25;
wire and26;
wire and27;
wire and28;
wire and29;
wire and30;
wire and31;
wire or3;
wire and32;
wire and33;
wire and34;
wire and35;
wire and36;
wire and37;
wire and38;
wire and39;
wire and40;
wire and41;
wire and42;
wire and43;
wire and44;
wire and45;
wire and46;
wire or4;

inv1$ in14_inv (.out(in14_not_weak), .in(in[14]));
inv1$ in13_inv (.out(in13_not_weak), .in(in[13]));
inv1$ in12_inv (.out(in12_not_weak), .in(in[12]));
inv1$ in11_inv (.out(in11_not_weak), .in(in[11]));
inv1$ in10_inv (.out(in10_not_weak), .in(in[10]));
inv1$ in9_inv (.out(in9_not_weak), .in(in[9]));
inv1$ in8_inv (.out(in8_not_weak), .in(in[8]));
inv1$ in7_inv (.out(in7_not_weak), .in(in[7]));
inv1$ in6_inv (.out(in6_not_weak), .in(in[6]));
inv1$ in5_inv (.out(in5_not_weak), .in(in[5]));
inv1$ in4_inv (.out(in4_not_weak), .in(in[4]));
inv1$ in3_inv (.out(in3_not_weak), .in(in[3]));
inv1$ in2_inv (.out(in2_not_weak), .in(in[2]));
inv1$ in1_inv (.out(in1_not_weak), .in(in[1]));
inv1$ in0_inv (.out(in0_not_weak), .in(in[0]));

bufferH16$ in14_buff(.out(in14_not), .in(in14_not_weak));
bufferH16$ in13_buff(.out(in13_not), .in(in13_not_weak));
bufferH16$ in12_buff(.out(in12_not), .in(in12_not_weak));
bufferH64$ in11_buff(.out(in11_not), .in(in11_not_weak));
bufferH64$ in10_buff(.out(in10_not), .in(in10_not_weak));
bufferH64$ in9_buff(.out(in9_not), .in(in9_not_weak));
bufferH64$ in8_buff(.out(in8_not), .in(in8_not_weak));
bufferH64$ in7_buff(.out(in7_not), .in(in7_not_weak));
bufferH64$ in6_buff(.out(in6_not), .in(in6_not_weak));
bufferH64$ in5_buff(.out(in5_not), .in(in5_not_weak));
bufferH64$ in4_buff(.out(in4_not), .in(in4_not_weak));
bufferH64$ in3_buff(.out(in3_not), .in(in3_not_weak));
bufferH64$ in2_buff(.out(in2_not), .in(in2_not_weak));
bufferH64$ in1_buff(.out(in1_not), .in(in1_not_weak));
bufferH64$ in0_buff(.out(in0_not), .in(in0_not_weak));

and16$ and_gate0(.out(and0), .in0(in[15]), .in1(in14_not), .in2(in13_not), .in3(in12_not), .in4(in11_not), .in5(in10_not), .in6(in9_not), .in7(in8_not), .in8(in7_not), .in9(in6_not), .in10(in5_not), .in11(in4_not), .in12(in3_not), .in13(in2_not), .in14(in1_not), .in15(in0_not));
and15$ and_gate1(.out(and1), .in0(in[14]), .in1(in13_not), .in2(in12_not), .in3(in11_not), .in4(in10_not), .in5(in9_not), .in6(in8_not), .in7(in7_not), .in8(in6_not), .in9(in5_not), .in10(in4_not), .in11(in3_not), .in12(in2_not), .in13(in1_not), .in14(in0_not));
and14$ and_gate2(.out(and2), .in0(in[13]), .in1(in12_not), .in2(in11_not), .in3(in10_not), .in4(in9_not), .in5(in8_not), .in6(in7_not), .in7(in6_not), .in8(in5_not), .in9(in4_not), .in10(in3_not), .in11(in2_not), .in12(in1_not), .in13(in0_not));
and13$ and_gate3(.out(and3), .in0(in[12]), .in1(in11_not), .in2(in10_not), .in3(in9_not), .in4(in8_not), .in5(in7_not), .in6(in6_not), .in7(in5_not), .in8(in4_not), .in9(in3_not), .in10(in2_not), .in11(in1_not), .in12(in0_not));
and11$ and_gate4(.out(and4), .in0(in[10]), .in1(in9_not), .in2(in8_not), .in3(in7_not), .in4(in6_not), .in5(in5_not), .in6(in4_not), .in7(in3_not), .in8(in2_not), .in9(in1_not), .in10(in0_not));
and12$ and_gate5(.out(and5), .in0(in[11]), .in1(in10_not), .in2(in9_not), .in3(in8_not), .in4(in7_not), .in5(in6_not), .in6(in5_not), .in7(in4_not), .in8(in3_not), .in9(in2_not), .in10(in1_not), .in11(in0_not));
and9$ and_gate6(.out(and6), .in0(in[8]), .in1(in7_not), .in2(in6_not), .in3(in5_not), .in4(in4_not), .in5(in3_not), .in6(in2_not), .in7(in1_not), .in8(in0_not));
and10$ and_gate7(.out(and7), .in0(in[9]), .in1(in8_not), .in2(in7_not), .in3(in6_not), .in4(in5_not), .in5(in4_not), .in6(in3_not), .in7(in2_not), .in8(in1_not), .in9(in0_not));
and16$ and_gate8(.out(and8), .in0(in[15]), .in1(in14_not), .in2(in13_not), .in3(in12_not), .in4(in11_not), .in5(in10_not), .in6(in9_not), .in7(in8_not), .in8(in7_not), .in9(in6_not), .in10(in5_not), .in11(in4_not), .in12(in3_not), .in13(in2_not), .in14(in1_not), .in15(in0_not));
and15$ and_gate9(.out(and9), .in0(in[14]), .in1(in13_not), .in2(in12_not), .in3(in11_not), .in4(in10_not), .in5(in9_not), .in6(in8_not), .in7(in7_not), .in8(in6_not), .in9(in5_not), .in10(in4_not), .in11(in3_not), .in12(in2_not), .in13(in1_not), .in14(in0_not));
and14$ and_gate10(.out(and10), .in0(in[13]), .in1(in12_not), .in2(in11_not), .in3(in10_not), .in4(in9_not), .in5(in8_not), .in6(in7_not), .in7(in6_not), .in8(in5_not), .in9(in4_not), .in10(in3_not), .in11(in2_not), .in12(in1_not), .in13(in0_not));
and13$ and_gate11(.out(and11), .in0(in[12]), .in1(in11_not), .in2(in10_not), .in3(in9_not), .in4(in8_not), .in5(in7_not), .in6(in6_not), .in7(in5_not), .in8(in4_not), .in9(in3_not), .in10(in2_not), .in11(in1_not), .in12(in0_not));
and7$ and_gate12(.out(and12), .in0(in[6]), .in1(in5_not), .in2(in4_not), .in3(in3_not), .in4(in2_not), .in5(in1_not), .in6(in0_not));
and6$ and_gate13(.out(and13), .in0(in[5]), .in1(in4_not), .in2(in3_not), .in3(in2_not), .in4(in1_not), .in5(in0_not));
and8$ and_gate14(.out(and14), .in0(in[7]), .in1(in6_not), .in2(in5_not), .in3(in4_not), .in4(in3_not), .in5(in2_not), .in6(in1_not), .in7(in0_not));
and5$ and_gate15(.out(and15), .in0(in[4]), .in1(in3_not), .in2(in2_not), .in3(in1_not), .in4(in0_not));
and16$ and_gate16(.out(and16), .in0(in[15]), .in1(in14_not), .in2(in13_not), .in3(in12_not), .in4(in11_not), .in5(in10_not), .in6(in9_not), .in7(in8_not), .in8(in7_not), .in9(in6_not), .in10(in5_not), .in11(in4_not), .in12(in3_not), .in13(in2_not), .in14(in1_not), .in15(in0_not));
and15$ and_gate17(.out(and17), .in0(in[14]), .in1(in13_not), .in2(in12_not), .in3(in11_not), .in4(in10_not), .in5(in9_not), .in6(in8_not), .in7(in7_not), .in8(in6_not), .in9(in5_not), .in10(in4_not), .in11(in3_not), .in12(in2_not), .in13(in1_not), .in14(in0_not));
and11$ and_gate18(.out(and18), .in0(in[10]), .in1(in9_not), .in2(in8_not), .in3(in7_not), .in4(in6_not), .in5(in5_not), .in6(in4_not), .in7(in3_not), .in8(in2_not), .in9(in1_not), .in10(in0_not));
and12$ and_gate19(.out(and19), .in0(in[11]), .in1(in10_not), .in2(in9_not), .in3(in8_not), .in4(in7_not), .in5(in6_not), .in6(in5_not), .in7(in4_not), .in8(in3_not), .in9(in2_not), .in10(in1_not), .in11(in0_not));
and7$ and_gate20(.out(and20), .in0(in[6]), .in1(in5_not), .in2(in4_not), .in3(in3_not), .in4(in2_not), .in5(in1_not), .in6(in0_not));
and4$ and_gate21(.out(and21), .in0(in[3]), .in1(in2_not), .in2(in1_not), .in3(in0_not));
and8$ and_gate22(.out(and22), .in0(in[7]), .in1(in6_not), .in2(in5_not), .in3(in4_not), .in4(in3_not), .in5(in2_not), .in6(in1_not), .in7(in0_not));
and3$ and_gate23(.out(and23), .in0(in[2]), .in1(in1_not), .in2(in0_not));
and16$ and_gate24(.out(and24), .in0(in[15]), .in1(in14_not), .in2(in13_not), .in3(in12_not), .in4(in11_not), .in5(in10_not), .in6(in9_not), .in7(in8_not), .in8(in7_not), .in9(in6_not), .in10(in5_not), .in11(in4_not), .in12(in3_not), .in13(in2_not), .in14(in1_not), .in15(in0_not));
and14$ and_gate25(.out(and25), .in0(in[13]), .in1(in12_not), .in2(in11_not), .in3(in10_not), .in4(in9_not), .in5(in8_not), .in6(in7_not), .in7(in6_not), .in8(in5_not), .in9(in4_not), .in10(in3_not), .in11(in2_not), .in12(in1_not), .in13(in0_not));
and12$ and_gate26(.out(and26), .in0(in[11]), .in1(in10_not), .in2(in9_not), .in3(in8_not), .in4(in7_not), .in5(in6_not), .in6(in5_not), .in7(in4_not), .in8(in3_not), .in9(in2_not), .in10(in1_not), .in11(in0_not));
and10$ and_gate27(.out(and27), .in0(in[9]), .in1(in8_not), .in2(in7_not), .in3(in6_not), .in4(in5_not), .in5(in4_not), .in6(in3_not), .in7(in2_not), .in8(in1_not), .in9(in0_not));
and6$ and_gate28(.out(and28), .in0(in[5]), .in1(in4_not), .in2(in3_not), .in3(in2_not), .in4(in1_not), .in5(in0_not));
and4$ and_gate29(.out(and29), .in0(in[3]), .in1(in2_not), .in2(in1_not), .in3(in0_not));
and8$ and_gate30(.out(and30), .in0(in[7]), .in1(in6_not), .in2(in5_not), .in3(in4_not), .in4(in3_not), .in5(in2_not), .in6(in1_not), .in7(in0_not));
and2$ and_gate31(.out(and31), .in0(in[1]), .in1(in0_not));
and16$ and_gate32(.out(and32), .in0(in[15]), .in1(in14_not), .in2(in13_not), .in3(in12_not), .in4(in11_not), .in5(in10_not), .in6(in9_not), .in7(in8_not), .in8(in7_not), .in9(in6_not), .in10(in5_not), .in11(in4_not), .in12(in3_not), .in13(in2_not), .in14(in1_not), .in15(in0_not));
and15$ and_gate33(.out(and33), .in0(in[14]), .in1(in13_not), .in2(in12_not), .in3(in11_not), .in4(in10_not), .in5(in9_not), .in6(in8_not), .in7(in7_not), .in8(in6_not), .in9(in5_not), .in10(in4_not), .in11(in3_not), .in12(in2_not), .in13(in1_not), .in14(in0_not));
and14$ and_gate34(.out(and34), .in0(in[13]), .in1(in12_not), .in2(in11_not), .in3(in10_not), .in4(in9_not), .in5(in8_not), .in6(in7_not), .in7(in6_not), .in8(in5_not), .in9(in4_not), .in10(in3_not), .in11(in2_not), .in12(in1_not), .in13(in0_not));
and13$ and_gate35(.out(and35), .in0(in[12]), .in1(in11_not), .in2(in10_not), .in3(in9_not), .in4(in8_not), .in5(in7_not), .in6(in6_not), .in7(in5_not), .in8(in4_not), .in9(in3_not), .in10(in2_not), .in11(in1_not), .in12(in0_not));
and11$ and_gate36(.out(and36), .in0(in[10]), .in1(in9_not), .in2(in8_not), .in3(in7_not), .in4(in6_not), .in5(in5_not), .in6(in4_not), .in7(in3_not), .in8(in2_not), .in9(in1_not), .in10(in0_not));
and12$ and_gate37(.out(and37), .in0(in[11]), .in1(in10_not), .in2(in9_not), .in3(in8_not), .in4(in7_not), .in5(in6_not), .in6(in5_not), .in7(in4_not), .in8(in3_not), .in9(in2_not), .in10(in1_not), .in11(in0_not));
and9$ and_gate38(.out(and38), .in0(in[8]), .in1(in7_not), .in2(in6_not), .in3(in5_not), .in4(in4_not), .in5(in3_not), .in6(in2_not), .in7(in1_not), .in8(in0_not));
and10$ and_gate39(.out(and39), .in0(in[9]), .in1(in8_not), .in2(in7_not), .in3(in6_not), .in4(in5_not), .in5(in4_not), .in6(in3_not), .in7(in2_not), .in8(in1_not), .in9(in0_not));
and7$ and_gate40(.out(and40), .in0(in[6]), .in1(in5_not), .in2(in4_not), .in3(in3_not), .in4(in2_not), .in5(in1_not), .in6(in0_not));
and6$ and_gate41(.out(and41), .in0(in[5]), .in1(in4_not), .in2(in3_not), .in3(in2_not), .in4(in1_not), .in5(in0_not));
and4$ and_gate42(.out(and42), .in0(in[3]), .in1(in2_not), .in2(in1_not), .in3(in0_not));
and8$ and_gate43(.out(and43), .in0(in[7]), .in1(in6_not), .in2(in5_not), .in3(in4_not), .in4(in3_not), .in5(in2_not), .in6(in1_not), .in7(in0_not));
and5$ and_gate44(.out(and44), .in0(in[4]), .in1(in3_not), .in2(in2_not), .in3(in1_not), .in4(in0_not));
and3$ and_gate45(.out(and45), .in0(in[2]), .in1(in1_not), .in2(in0_not));
and2$ and_gate46(.out(and46), .in0(in[1]), .in1(in0_not));

or8$ or_gate0(.out(or0), .in0(and0), .in1(and1), .in2(and2), .in3(and3), .in4(and4), .in5(and5), .in6(and6), .in7(and7));
or8$ or_gate1(.out(or1), .in0(and8), .in1(and9), .in2(and10), .in3(and11), .in4(and12), .in5(and13), .in6(and14), .in7(and15));
or8$ or_gate2(.out(or2), .in0(and16), .in1(and17), .in2(and18), .in3(and19), .in4(and20), .in5(and21), .in6(and22), .in7(and23));
or8$ or_gate3(.out(or3), .in0(and24), .in1(and25), .in2(and26), .in3(and27), .in4(and28), .in5(and29), .in6(and30), .in7(and31));
or16$ or_gate4(.out(or4), .in0(and32), .in1(and33), .in2(and34), .in3(and35), .in4(and36), .in5(and37), .in6(and38), .in7(and39), .in8(and40), .in9(and41), .in10(and42), .in11(and43), .in12(and44), .in13(in[0]), .in14(and45), .in15(and46));

assign out[3] = or0;
assign out[2] = or1;
assign out[1] = or2;
assign out[0] = or3;
assign v = or4;

assign out[31:4] = 28'h0000000;

endmodule