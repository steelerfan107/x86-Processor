module opcode_modrm_control_cloud (
 input  sizeov,				    
 input 	modrm7, 
 input 	modrm6, 
 input 	modrm5, 
 input 	modrm4, 
 input 	modrm3, 
 input 	modrm2, 
 input 	modrm1, 
 input 	modrm0, 
 input 	op15, 
 input 	op14, 
 input 	op13, 
 input 	op12, 
 input 	op11, 
 input 	op10, 
 input 	op9, 
 input 	op8, 
 input 	op7, 
 input 	op6, 
 input 	op5, 
 input 	op4, 
 input 	op3, 
 input 	op2, 
 input 	op1, 
 input 	op0,
 output setd, 
 output cleard, 
 output size2, 
 output size1, 
 output size0, 
 output op0_2, 
 output op0_1, 
 output op0_0, 
 output op1_2, 
 output op1_1, 
 output op1_0, 
 output op0_reg_4, 
 output op0_reg_3, 
 output op0_reg_2, 
 output op0_reg_1, 
 output op0_reg_0, 
 output op1_reg_4, 
 output op1_reg_3, 
 output op1_reg_2, 
 output op1_reg_1, 
 output op1_reg_0, 
 output alu_op_3, 
 output alu_op_2, 
 output alu_op_1, 
 output alu_op_0, 
 output flag0_2, 
 output flag0_1, 
 output flag0_0, 
 output flag1_2, 
 output flag1_1, 
 output flag1_0, 
 output stack_op_1, 
 output stack_op_0, 
 output rom_control_2, 
 output rom_control_1, 
 output rom_control_0				   
);

wire sizeov_not;
wire modrm7_not;
wire modrm6_not;
wire modrm5_not;
wire modrm2_not;
wire modrm0_not;
wire op15_not;
wire op14_not;
wire op13_not;
wire op12_not;
wire op11_not;
wire op10_not;
wire op9_not;
wire op8_not;
wire op7_not;
wire op6_not;
wire op5_not;
wire op2_not;
wire op1_not;
wire and0;
wire modrm4_not;
wire modrm1_not;
wire and1;
wire op5_not;
wire op4_not;
wire and2;
wire modrm3_not;
wire op14_not;
wire op3_not;
wire and3;
wire sizeov_not;
wire and4;
wire and5;
wire sizeov_not;
wire op15_not;
wire and6;
wire op2_not;
wire and7;
wire modrm0_not;
wire and8;
wire modrm3_not;
wire and9;
wire modrm6_not;
wire and10;
wire modrm1_not;
wire and11;
wire and12;
wire and13;
wire or0;
wire and14;
wire and15;
wire modrm1_not;
wire and16;
wire and17;
wire op12_not;
wire and18;
wire and19;
wire modrm5_not;
wire and20;
wire and21;
wire and22;
wire op11_not;
wire and23;
wire op10_not;
wire and24;
wire and25;
wire or1;
wire and26;
wire op7_not;
wire and27;
wire modrm2_not;
wire and28;
wire modrm0_not;
wire and29;
wire and30;
wire and31;
wire and32;
wire and33;
wire and34;
wire and35;
wire modrm7_not;
wire and36;
wire and37;
wire and38;
wire and39;
wire or2;
wire and40;
wire and41;
wire and42;
wire and43;
wire modrm4_not;
wire and44;
wire and45;
wire modrm7_not;
wire and46;
wire modrm5_not;
wire and47;
wire or3;
wire and48;
wire and49;
wire and50;
wire and51;
wire and52;
wire and53;
wire and54;
wire and55;
wire and56;
wire and57;
wire and58;
wire and59;
wire and60;
wire and61;
wire or4;
wire and62;
wire and63;
wire and64;
wire and65;
wire and66;
wire and67;
wire and68;
wire and69;
wire and70;
wire and71;
wire and72;
wire and73;
wire and74;
wire and75;
wire and76;
wire and77;
wire and78;
wire and79;
wire or5;
wire and80;
wire and81;
wire and82;
wire and83;
wire and84;
wire and85;
wire and86;
wire op6_not;
wire and87;
wire and88;
wire op3_not;
wire and89;
wire and90;
wire modrm3_not;
wire and91;
wire and92;
wire and93;
wire modrm6_not;
wire and94;
wire and95;
wire modrm4_not;
wire and96;
wire and97;
wire and98;
wire or6;
wire and99;
wire and100;
wire and101;
wire op4_not;
wire and102;
wire and103;
wire and104;
wire and105;
wire and106;
wire and107;
wire and108;
wire and109;
wire and110;
wire and111;
wire and112;
wire and113;
wire and114;
wire and115;
wire or7;
wire and116;
wire and117;
wire and118;
wire and119;
wire op9_not;
wire and120;
wire and121;
wire and122;
wire and123;
wire and124;
wire and125;
wire and126;
wire and127;
wire op8_not;
wire and128;
wire and129;
wire and130;
wire and131;
wire or8;
wire and132;
wire and133;
wire and134;
wire and135;
wire and136;
wire and137;
wire and138;
wire and139;
wire and140;
wire and141;
wire and142;
wire and143;
wire op15_not;
wire and144;
wire and145;
wire or9;
wire and146;
wire and147;
wire and148;
wire and149;
wire and150;
wire and151;
wire and152;
wire and153;
wire and154;
wire and155;
wire and156;
wire and157;
wire and158;
wire and159;
wire and160;
wire and161;
wire and162;
wire and163;
wire op14_not;
wire and164;
wire or10;
wire and165;
wire and166;
wire and167;
wire and168;
wire and169;
wire and170;
wire op13_not;
wire and171;
wire and172;
wire and173;
wire and174;
wire and175;
wire and176;
wire and177;
wire and178;
wire and179;
wire and180;
wire and181;
wire and182;
wire and183;
wire and184;
wire and185;
wire and186;
wire and187;
wire and188;
wire or11;
wire and189;
wire and190;
wire and191;
wire and192;
wire and193;
wire and194;
wire and195;
wire and196;
wire and197;
wire and198;
wire and199;
wire and200;
wire and201;
wire and202;
wire and203;
wire and204;
wire and205;
wire and206;
wire and207;
wire and208;
wire and209;
wire and210;
wire and211;
wire and212;
wire and213;
wire and214;
wire or12;
wire and215;
wire and216;
wire and217;
wire and218;
wire and219;
wire and220;
wire and221;
wire and222;
wire and223;
wire and224;
wire and225;
wire and226;
wire and227;
wire and228;
wire and229;
wire and230;
wire and231;
wire and232;
wire and233;
wire and234;
wire and235;
wire and236;
wire and237;
wire and238;
wire or13;
wire and239;
wire and240;
wire and241;
wire and242;
wire and243;
wire and244;
wire and245;
wire and246;
wire and247;
wire and248;
wire and249;
wire and250;
wire and251;
wire and252;
wire and253;
wire and254;
wire and255;
wire and256;
wire and257;
wire and258;
wire and259;
wire and260;
wire and261;
wire or14;
wire and262;
wire and263;
wire and264;
wire and265;
wire and266;
wire and267;
wire and268;
wire and269;
wire and270;
wire and271;
wire and272;
wire and273;
wire and274;
wire and275;
wire and276;
wire and277;
wire and278;
wire and279;
wire and280;
wire and281;
wire or15;
wire and282;
wire and283;
wire and284;
wire and285;
wire and286;
wire and287;
wire and288;
wire and289;
wire and290;
wire and291;
wire and292;
wire and293;
wire and294;
wire and295;
wire and296;
wire and297;
wire or16;
wire and298;
wire and299;
wire and300;
wire and301;
wire and302;
wire and303;
wire and304;
wire and305;
wire and306;
wire and307;
wire and308;
wire and309;
wire and310;
wire and311;
wire and312;
wire and313;
wire and314;
wire and315;
wire and316;
wire and317;
wire and318;
wire and319;
wire or17;
wire and320;
wire and321;
wire and322;
wire and323;
wire and324;
wire and325;
wire and326;
wire and327;
wire and328;
wire and329;
wire and330;
wire and331;
wire and332;
wire and333;
wire and334;
wire and335;
wire and336;
wire and337;
wire and338;
wire or18;
wire and339;
wire and340;
wire and341;
wire and342;
wire and343;
wire and344;
wire and345;
wire and346;
wire and347;
wire and348;
wire and349;
wire and350;
wire and351;
wire and352;
wire and353;
wire and354;
wire and355;
wire or19;
wire and356;
wire and357;
wire and358;
wire and359;
wire and360;
wire and361;
wire and362;
wire and363;
wire and364;
wire and365;
wire and366;
wire and367;
wire and368;
wire and369;
wire and370;
wire and371;
wire and372;
wire and373;
wire and374;
wire or20;
wire and375;
wire and376;
wire and377;
wire and378;
wire and379;
wire and380;
wire and381;
wire and382;
wire and383;
wire and384;
wire and385;
wire and386;
wire and387;
wire and388;
wire and389;
wire and390;
wire and391;
wire or21;
wire and392;
wire and393;
wire and394;
wire and395;
wire and396;
wire and397;
wire and398;
wire and399;
wire and400;
wire and401;
wire and402;
wire and403;
wire and404;
wire and405;
wire and406;
wire and407;
wire and408;
wire and409;
wire and410;
wire or22;
wire and411;
wire and412;
wire and413;
wire and414;
wire and415;
wire and416;
wire and417;
wire and418;
wire and419;
wire and420;
wire and421;
wire and422;
wire or23;
wire and423;
wire and424;
wire and425;
wire and426;
wire and427;
wire and428;
wire and429;
wire and430;
wire and431;
wire and432;
wire and433;
wire and434;
wire or24;
wire and435;
wire and436;
wire and437;
wire and438;
wire and439;
wire and440;
wire and441;
wire and442;
wire and443;
wire and444;
wire and445;
wire and446;
wire or25;
wire and447;
wire and448;
wire and449;
wire and450;
wire and451;
wire and452;
wire and453;
wire and454;
wire and455;
wire and456;
wire or26;
wire and457;
wire and458;
wire and459;
wire and460;
wire and461;
wire and462;
wire and463;
wire and464;
wire and465;
wire and466;
wire modrm2_not;
wire and467;
wire and468;
wire and469;
wire and470;
wire or27;
wire and471;
wire and472;
wire and473;
wire and474;
wire and475;
wire and476;
wire and477;
wire and478;
wire and479;
wire and480;
wire and481;
wire and482;
wire and483;
wire and484;
wire and485;
wire and486;
wire and487;
wire and488;
wire or28;
wire and489;
wire and490;
wire and491;
wire and492;
wire and493;
wire and494;
wire and495;
wire and496;
wire and497;
wire and498;
wire and499;
wire and500;
wire and501;
wire and502;
wire and503;
wire or29;
wire and504;
wire and505;
wire and506;
wire and507;
wire and508;
wire and509;
wire and510;
wire and511;
wire and512;
wire and513;
wire or30;
wire and514;
wire and515;
wire and516;
wire and517;
wire and518;
wire and519;
wire and520;
wire and521;
wire and522;
wire and523;
wire and524;
wire or31;
wire and525;
wire and526;
wire and527;
wire and528;
wire and529;
wire and530;
wire and531;
wire and532;
wire and533;
wire and534;
wire and535;
wire or32;
wire and536;
wire and537;
wire and538;
wire and539;
wire and540;
wire and541;
wire and542;
wire and543;
wire and544;
wire and545;
wire and546;
wire and547;
wire and548;
wire or33;
wire and549;
wire and550;
wire and551;
wire and552;
wire and553;
wire and554;
wire and555;
wire and556;
wire and557;
wire and558;
wire and559;
wire and560;
wire and561;
wire and562;
wire and563;
wire or34;
wire and564;
wire and565;
wire and566;
wire and567;
wire and568;
wire and569;
wire and570;
wire and571;
wire and572;
wire and573;
wire and574;
wire and575;
wire and576;
wire and577;
wire or35;

inv1$ sizeov_inv (.out(sizeov_not), .in(sizeov));
inv1$ modrm7_inv (.out(modrm7_not), .in(modrm7));
inv1$ modrm6_inv (.out(modrm6_not), .in(modrm6));
inv1$ modrm5_inv (.out(modrm5_not), .in(modrm5));
inv1$ modrm2_inv (.out(modrm2_not), .in(modrm2));
inv1$ modrm0_inv (.out(modrm0_not), .in(modrm0));
inv1$ op15_inv (.out(op15_not), .in(op15));
inv1$ op14_inv (.out(op14_not), .in(op14));
inv1$ op13_inv (.out(op13_not), .in(op13));
inv1$ op12_inv (.out(op12_not), .in(op12));
inv1$ op11_inv (.out(op11_not), .in(op11));
inv1$ op10_inv (.out(op10_not), .in(op10));
inv1$ op9_inv (.out(op9_not), .in(op9));
inv1$ op8_inv (.out(op8_not), .in(op8));
inv1$ op7_inv (.out(op7_not), .in(op7));
inv1$ op6_inv (.out(op6_not), .in(op6));
inv1$ op5_inv (.out(op5_not), .in(op5));
inv1$ op2_inv (.out(op2_not), .in(op2));
inv1$ op1_inv (.out(op1_not), .in(op1));
inv1$ modrm4_inv (.out(modrm4_not), .in(modrm4));
inv1$ modrm1_inv (.out(modrm1_not), .in(modrm1));
inv1$ op5_inv (.out(op5_not), .in(op5));
inv1$ op4_inv (.out(op4_not), .in(op4));
inv1$ modrm3_inv (.out(modrm3_not), .in(modrm3));
inv1$ op14_inv (.out(op14_not), .in(op14));
inv1$ op3_inv (.out(op3_not), .in(op3));
inv1$ sizeov_inv (.out(sizeov_not), .in(sizeov));
inv1$ sizeov_inv (.out(sizeov_not), .in(sizeov));
inv1$ op15_inv (.out(op15_not), .in(op15));
inv1$ op2_inv (.out(op2_not), .in(op2));
inv1$ modrm0_inv (.out(modrm0_not), .in(modrm0));
inv1$ modrm3_inv (.out(modrm3_not), .in(modrm3));
inv1$ modrm6_inv (.out(modrm6_not), .in(modrm6));
inv1$ modrm1_inv (.out(modrm1_not), .in(modrm1));
inv1$ modrm1_inv (.out(modrm1_not), .in(modrm1));
inv1$ op12_inv (.out(op12_not), .in(op12));
inv1$ modrm5_inv (.out(modrm5_not), .in(modrm5));
inv1$ op11_inv (.out(op11_not), .in(op11));
inv1$ op10_inv (.out(op10_not), .in(op10));
inv1$ op7_inv (.out(op7_not), .in(op7));
inv1$ modrm2_inv (.out(modrm2_not), .in(modrm2));
inv1$ modrm0_inv (.out(modrm0_not), .in(modrm0));
inv1$ modrm7_inv (.out(modrm7_not), .in(modrm7));
inv1$ modrm4_inv (.out(modrm4_not), .in(modrm4));
inv1$ modrm7_inv (.out(modrm7_not), .in(modrm7));
inv1$ modrm5_inv (.out(modrm5_not), .in(modrm5));
inv1$ op6_inv (.out(op6_not), .in(op6));
inv1$ op3_inv (.out(op3_not), .in(op3));
inv1$ modrm3_inv (.out(modrm3_not), .in(modrm3));
inv1$ modrm6_inv (.out(modrm6_not), .in(modrm6));
inv1$ modrm4_inv (.out(modrm4_not), .in(modrm4));
inv1$ op4_inv (.out(op4_not), .in(op4));
inv1$ op9_inv (.out(op9_not), .in(op9));
inv1$ op8_inv (.out(op8_not), .in(op8));
inv1$ op15_inv (.out(op15_not), .in(op15));
inv1$ op14_inv (.out(op14_not), .in(op14));
inv1$ op13_inv (.out(op13_not), .in(op13));
inv1$ modrm2_inv (.out(modrm2_not), .in(modrm2));

and24$ and_gate0(.out(and0), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3), .in6(modrm2_not), .in7(modrm1
), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not), .in19(op5_not), .in20(op4), .in21(op3), .in22(op2_not), .in23(op1_not));
and20$ and_gate1(.out(and1), .in0(modrm4_not), .in1(modrm3), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0_not), .in5(op15
), .in6(op14_not), .in7(op13_not), .in8(op12_not), .in9(op11_not), .in10(op10_not), .in11(op9), .in12(op8), .in13(op7_not), .in14(op6), .in15(op5), .in16(op4), .in17(op3), .in18(op2), .in19(op1));
and16$ and_gate2(.out(and2), .in0(
sizeov), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(modrm4), .in5(modrm3), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6
), .in11(op5_not), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1_not));
and19$ and_gate3(.out(and3), .in0(modrm3_not), .in1(modrm2_not), .in2(modrm1_not), .in3(modrm0_not), .in4(op15), .in5(op14_not), .in6(op13), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8_not), .in12(op7_not), .in13(op6_not), .in14(op5_not), .in15(op4_not), .in16(op3_not), .in17(op2_not), .in18(op1_not));
and16$ and_gate4(.out(and4), .in0(sizeov_not), .in1(modrm7), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4
), .in13(op3_not), .in14(op2), .in15(op1_not));
and18$ and_gate5(.out(and5), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11
), .in8(op10_not), .in9(op9_not), .in10(op8_not), .in11(op7_not), .in12(op6_not), .in13(op5_not), .in14(op4_not), .in15(op3_not), .in16(op2_not), .in17(op1_not));
and16$ and_gate6(.out(and6), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3), .in6(modrm2_not), .in7(modrm1), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12), .in13(op6_not), .in14(op5), .in15(op1));
and16$ and_gate7(.out(and7), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5
), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15), .in10(op14), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1));
and15$ and_gate8(.out(and8), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15_not), .in9(op14_not), .in10(op13), .in11(op7_not), .in12(op6), .in13(op2), .in14(op1));
and14$ and_gate9(.out(and9), .in0(modrm6), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(modrm2_not), .in5(modrm1_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3), .in12(op2), .in13(op1));
and16$ and_gate10(.out(and10), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and13$ and_gate11(.out(and11), .in0(modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(modrm1_not), .in5(modrm0), .in6(op7_not), .in7(op6_not), .in8(op5_not), .in9(op4_not), .in10(op3), .in11(op2), .in12(op1));
and10$ and_gate12(.out(and12), .in0(modrm2_not), .in1(modrm1), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13), .in6(op4_not), .in7(op3), .in8(op2), .in9(op1_not));
and10$ and_gate13(.out(and13), .in0(sizeov), .in1(modrm7_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11), .in8(op2_not), .in9(op1_not));
and23$ and_gate14(.out(and14), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5), .in4(modrm4), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6), .in19(op5_not), .in20(op4_not), .in21(op3_not), .in22(op1));
and20$ and_gate15(.out(and15), .in0(modrm4_not), .in1(modrm3), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0_not), .in5(op15), .in6(op14_not), .in7(op13_not), .in8(op12_not), .in9(op11_not), .in10(op10_not), .in11(op9), .in12(op8), .in13(op7_not), .in14(op6), .in15(op5), .in16(op4), .in17(op3), .in18(op2), .in19(op1));
and17$ and_gate16(.out(and16), .in0(modrm1_not), .in1(modrm0_not), .in2(op15_not), .in3(op14_not), .in4(op13), .in5(op12), .in6(op11), .in7(op10), .in8(op9), .in9(op8), .in10(op7), .in11(op6), .in12(op5
), .in13(op4), .in14(op3_not), .in15(op2), .in16(op1_not));
and20$ and_gate17(.out(and17), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13_not), .in8(op12_not), .in9(op11_not), .in10(op10_not), .in11(op9), .in12(op8_not), .in13(op7_not), .in14(op6), .in15(op5_not), .in16(op4_not), .in17(op3_not), .in18(op2_not), .in19(op1_not));
and19$ and_gate18(.out(and18), .in0(modrm3_not), .in1(modrm2_not), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8), .in12(op7_not), .in13(op6_not), .in14(op5), .in15(op4_not), .in16(op3_not), .in17(op2_not), .in18(op1_not));
and16$ and_gate19(.out(and19), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3), .in6(modrm2_not), .in7(modrm1), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12), .in13(op6_not), .in14(op5), .in15(op1));
and16$ and_gate20(.out(and20), .in0(sizeov), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4), .in13(op3_not), .in14(op2
), .in15(op1_not));
and13$ and_gate21(.out(and21), .in0(modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(modrm1_not), .in5(modrm0), .in6(op7_not), .in7(op6_not), .in8(op5_not), .in9(op4_not), .in10(op3), .in11(op2), .in12(op1));
and10$ and_gate22(.out(and22), .in0(sizeov_not), .in1(modrm1_not), .in2(modrm0), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op3_not), .in8(op2), .in9(op1));
and10$ and_gate23(.out(and23), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op1_not));
and10$ and_gate24(.out(and24), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and8$ and_gate25(.out(and25), .in0(op14), .in1(op13), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and24$ and_gate26(.out(and26), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3), .in6(modrm2_not), .in7(modrm1
), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not), .in19(op5_not), .in20(op4), .in21(op3), .in22(op2_not), .in23(op1_not));
and20$ and_gate27(.out(and27), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3
), .in6(modrm2), .in7(modrm1), .in8(modrm0), .in9(op15_not), .in10(op14_not), .in11(op13), .in12(op12_not), .in13(op11), .in14(op10), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6), .in19(op5));
and18$ and_gate28(.out(and28), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9), .in16(op3_not), .in17(op2));
and16$ and_gate29(.out(and29), .in0(modrm0_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4), .in13(op3
), .in14(op2), .in15(op1_not));
and16$ and_gate30(.out(and30), .in0(sizeov_not), .in1(modrm7), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3), .in14(op2_not), .in15(op1));
and19$ and_gate31(.out(and31), .in0(modrm3_not), .in1(modrm2_not), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8), .in12(op7_not), .in13(op6_not), .in14(op5), .in15(op4_not), .in16(op3_not), .in17(op2_not), .in18(op1_not));
and18$ and_gate32(.out(and32), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14
), .in5(op13_not), .in6(op12), .in7(op11), .in8(op10_not), .in9(op9_not), .in10(op8_not), .in11(op7_not), .in12(op6_not), .in13(op5_not), .in14(op4_not), .in15(op3_not), .in16(op2_not), .in17(op1_not));
and14$ and_gate33(.out(and33), .in0(
modrm6), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(modrm2_not), .in5(modrm1_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3), .in12(op2), .in13(op1));
and16$ and_gate34(.out(and34), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and10$ and_gate35(.out(and35), .in0(modrm2_not), .in1(modrm1
), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13), .in6(op4_not), .in7(op3), .in8(op2), .in9(op1_not));
and10$ and_gate36(.out(and36), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm0_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op2_not), .in9(op1_not));
and10$ and_gate37(.out(and37), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op15_not), .in4(op14), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op1_not));
and10$ and_gate38(.out(and38), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate39(.out(and39), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not));
and17$ and_gate40(.out(and40), .in0(modrm1_not), .in1(modrm0_not), .in2(op15_not), .in3(op14_not), .in4(op13), .in5(op12), .in6(op11), .in7(op10), .in8(op9), .in9(op8), .in10(op7), .in11(op6
), .in12(op5), .in13(op4), .in14(op3_not), .in15(op2), .in16(op1_not));
and16$ and_gate41(.out(and41), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10
), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1));
and16$ and_gate42(.out(and42), .in0(sizeov), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4
), .in13(op3_not), .in14(op2), .in15(op1_not));
and16$ and_gate43(.out(and43), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and13$ and_gate44(.out(and44), .in0(modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(modrm1_not), .in5(modrm0), .in6(op7_not), .in7(op6_not), .in8(op5_not), .in9(op4_not), .in10(op3), .in11(op2), .in12(op1));
and10$ and_gate45(.out(and45), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm0_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op2_not), .in9(op1_not));
and10$ and_gate46(.out(and46), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate47(.out(and47), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not));
and19$ and_gate48(.out(and48), .in0(modrm3_not), .in1(modrm2_not), .in2(modrm1_not), .in3(modrm0_not), .in4(op15), .in5(op14_not), .in6(op13), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8_not), .in12(op7_not), .in13(op6_not), .in14(op5_not), .in15(op4_not), .in16(op3_not), .in17(op2_not), .in18(op1_not));
and16$ and_gate49(.out(and49), .in0(modrm0_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not));
and16$ and_gate50(.out(and50), .in0(sizeov_not), .in1(modrm7), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3), .in14(op2_not), .in15(op1));
and18$ and_gate51(.out(and51), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11), .in8(op10_not), .in9(op9_not), .in10(op8_not), .in11(op7_not), .in12(op6_not), .in13(op5_not), .in14(op4_not), .in15(op3_not), .in16(op2_not), .in17(op1_not));
and17$ and_gate52(.out(and52), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8));
and16$ and_gate53(.out(and53), .in0(
sizeov), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate54(.out(and54), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and10$ and_gate55(.out(and55), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not));
and10$ and_gate56(.out(and56), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm0_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op2_not), .in9(op1_not));
and10$ and_gate57(.out(and57), .in0(sizeov
), .in1(modrm7_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11), .in8(op2_not), .in9(op1_not));
and10$ and_gate58(.out(and58), .in0(sizeov_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op3_not), .in8(op2_not), .in9(op1));
and10$ and_gate59(.out(and59), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op15_not), .in4(op14), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op1_not));
and10$ and_gate60(.out(and60), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not));
and10$ and_gate61(.out(and61), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and17$ and_gate62(.out(and62), .in0(modrm1_not), .in1(modrm0_not), .in2(op15_not), .in3(op14_not), .in4(op13), .in5(op12), .in6(op11), .in7(op10), .in8(op9), .in9(op8), .in10(op7), .in11(op6
), .in12(op5), .in13(op4), .in14(op3_not), .in15(op2), .in16(op1_not));
and19$ and_gate63(.out(and63), .in0(modrm3_not), .in1(modrm2_not), .in2(modrm1_not), .in3(modrm0_not), .in4(op15), .in5(op14_not), .in6(op13), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8_not), .in12(op7_not), .in13(op6_not), .in14(op5_not), .in15(op4_not), .in16(op3_not), .in17(op2_not), .in18(op1_not));
and16$ and_gate64(.out(and64), .in0(sizeov_not), .in1(modrm7), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4
), .in13(op3_not), .in14(op2), .in15(op1_not));
and16$ and_gate65(.out(and65), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8
), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1));
and18$ and_gate66(.out(and66), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14
), .in5(op13_not), .in6(op12), .in7(op11), .in8(op10_not), .in9(op9_not), .in10(op8_not), .in11(op7_not), .in12(op6_not), .in13(op5_not), .in14(op4_not), .in15(op3_not), .in16(op2_not), .in17(op1_not));
and16$ and_gate67(.out(and67), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15), .in10(op14), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1));
and16$ and_gate68(.out(and68), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and13$ and_gate69(.out(and69), .in0(
modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(modrm1_not), .in5(modrm0), .in6(op7_not), .in7(op6_not), .in8(op5_not), .in9(op4_not), .in10(op3
), .in11(op2), .in12(op1));
and10$ and_gate70(.out(and70), .in0(modrm3_not), .in1(modrm2), .in2(modrm1), .in3(modrm0_not), .in4(op9_not), .in5(op8_not), .in6(op7), .in7(op6_not), .in8(op5_not), .in9(op4_not));
and10$ and_gate71(.out(and71), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not));
and10$ and_gate72(.out(and72), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op14_not), .in5(op13), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate73(.out(and73), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op15_not), .in4(op14), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op1_not));
and10$ and_gate74(.out(and74), .in0(
modrm0), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op6_not), .in5(op5_not), .in6(op4_not), .in7(op3_not), .in8(op2_not), .in9(op1_not));
and10$ and_gate75(.out(and75), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op1_not));
and10$ and_gate76(.out(and76), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate77(.out(and77), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8_not));
and10$ and_gate78(.out(and78), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not));
and10$ and_gate79(.out(and79), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and19$ and_gate80(.out(and80), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9), .in16(op8), .in17(op7), .in18(op6));
and17$ and_gate81(.out(and81), .in0(modrm1_not), .in1(modrm0_not), .in2(op15_not), .in3(op14_not), .in4(op13), .in5(op12), .in6(op11), .in7(op10), .in8(op9), .in9(op8), .in10(op7), .in11(op6), .in12(op5
), .in13(op4), .in14(op3_not), .in15(op2), .in16(op1_not));
and16$ and_gate82(.out(and82), .in0(modrm0_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10), .in7(op9
), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not));
and18$ and_gate83(.out(and83), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8), .in17(op7));
and18$ and_gate84(.out(and84), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14), .in5(op13_not), .in6(op12
), .in7(op11), .in8(op10_not), .in9(op9_not), .in10(op8_not), .in11(op7_not), .in12(op6_not), .in13(op5_not), .in14(op4_not), .in15(op3_not), .in16(op2_not), .in17(op1_not));
and17$ and_gate85(.out(and85), .in0(sizeov
), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15
), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8));
and16$ and_gate86(.out(and86), .in0(sizeov_not), .in1(modrm7_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op8_not), .in9(op7), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate87(.out(and87), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate88(.out(and88), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and14$ and_gate89(.out(and89), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0), .in5(op15), .in6(op14), .in7(op13_not), .in8(op12_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and10$ and_gate90(.out(and90), .in0(modrm2_not), .in1(modrm1), .in2(modrm0), .in3(op15_not), .in4(op8), .in5(op7_not), .in6(op6), .in7(op5_not), .in8(op4), .in9(op3_not));
and10$ and_gate91(.out(and91), .in0(modrm3_not), .in1(modrm2), .in2(modrm1), .in3(modrm0_not), .in4(op9_not), .in5(op8_not), .in6(op7), .in7(op6_not), .in8(op5_not), .in9(op4_not));
and10$ and_gate92(.out(and92), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op14_not), .in5(op13), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate93(.out(and93), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op1_not));
and10$ and_gate94(.out(and94), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not));
and10$ and_gate95(.out(and95), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8_not));
and10$ and_gate96(.out(and96), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not));
and10$ and_gate97(.out(and97), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate98(.out(and98), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not));
and17$ and_gate99(.out(and99), .in0(modrm1_not), .in1(modrm0_not), .in2(op15_not), .in3(op14_not), .in4(op13), .in5(op12), .in6(op11), .in7(op10), .in8(op9), .in9(op8), .in10(op7), .in11(op6
), .in12(op5), .in13(op4), .in14(op3_not), .in15(op2), .in16(op1_not));
and16$ and_gate100(.out(and100), .in0(sizeov_not), .in1(modrm7), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4), .in13(op3_not), .in14(op2), .in15(op1_not));
and16$ and_gate101(.out(and101), .in0(modrm0_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not));
and16$ and_gate102(.out(and102), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1));
and18$ and_gate103(.out(and103), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8
), .in17(op7));
and16$ and_gate104(.out(and104), .in0(sizeov_not), .in1(modrm7_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op8_not), .in9(op7
), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and14$ and_gate105(.out(and105), .in0(modrm6), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(modrm2_not), .in5(modrm1_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3), .in12(op2), .in13(op1));
and16$ and_gate106(.out(and106), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and10$ and_gate107(.out(and107), .in0(modrm2_not), .in1(modrm1), .in2(modrm0), .in3(op15_not), .in4(op8), .in5(op7_not), .in6(op6), .in7(op5_not), .in8(op4), .in9(op3_not));
and10$ and_gate108(.out(and108), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3), .in6(op8), .in7(op7
), .in8(op6_not), .in9(op5));
and10$ and_gate109(.out(and109), .in0(modrm1_not), .in1(modrm0), .in2(op15), .in3(op14_not), .in4(op7), .in5(op6_not), .in6(op5), .in7(op4_not), .in8(op3), .in9(op2_not));
and10$ and_gate110(.out(and110), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not));
and10$ and_gate111(.out(and111), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8_not));
and10$ and_gate112(.out(and112), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not));
and10$ and_gate113(.out(and113), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate114(.out(and114), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not));
and8$ and_gate115(.out(and115), .in0(
op14), .in1(op13), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and16$ and_gate116(.out(and116), .in0(modrm0_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4
), .in13(op3), .in14(op2), .in15(op1_not));
and16$ and_gate117(.out(and117), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8
), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1));
and16$ and_gate118(.out(and118), .in0(sizeov), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate119(.out(and119), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate120(.out(and120), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate121(.out(and121), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate122(.out(and122), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and13$ and_gate123(.out(and123), .in0(modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(modrm1_not), .in5(modrm0), .in6(op7_not), .in7(op6_not), .in8(op5_not), .in9(op4_not), .in10(op3), .in11(op2), .in12(op1));
and10$ and_gate124(.out(and124), .in0(modrm1_not), .in1(modrm0), .in2(op15), .in3(op14_not), .in4(op7), .in5(op6_not), .in6(op5), .in7(op4_not), .in8(op3), .in9(op2_not));
and10$ and_gate125(.out(and125), .in0(modrm0), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op6_not), .in5(op5_not), .in6(op4_not), .in7(op3_not), .in8(op2_not), .in9(op1_not));
and10$ and_gate126(.out(and126), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not));
and10$ and_gate127(.out(and127), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8_not));
and10$ and_gate128(.out(and128), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not));
and10$ and_gate129(.out(and129), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate130(.out(and130), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not));
and8$ and_gate131(.out(and131), .in0(sizeov), .in1(op13), .in2(op12), .in3(op11_not), .in4(op10_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and19$ and_gate132(.out(and132), .in0(modrm3_not), .in1(modrm2_not), .in2(modrm1_not), .in3(modrm0_not), .in4(op15), .in5(op14_not), .in6(op13), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8_not), .in12(op7_not), .in13(op6_not), .in14(op5_not), .in15(op4_not), .in16(op3_not), .in17(op2_not), .in18(op1_not));
and16$ and_gate133(.out(and133), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1));
and17$ and_gate134(.out(and134), .in0(
sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8));
and16$ and_gate135(.out(and135), .in0(sizeov), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate136(.out(and136), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and14$ and_gate137(.out(and137), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0
), .in5(op15), .in6(op14), .in7(op13_not), .in8(op12_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and13$ and_gate138(.out(and138), .in0(sizeov_not), .in1(modrm7
), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op12), .in8(op11), .in9(op10_not), .in10(op9_not), .in11(op2_not), .in12(op1_not));
and13$ and_gate139(.out(and139), .in0(modrm3_not), .in1(modrm2), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not));
and10$ and_gate140(.out(and140), .in0(modrm3_not), .in1(modrm2), .in2(modrm1), .in3(modrm0_not), .in4(op9_not), .in5(op8_not), .in6(op7), .in7(op6_not), .in8(op5_not), .in9(op4_not));
and10$ and_gate141(.out(and141), .in0(modrm0), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op6_not), .in5(op5_not), .in6(op4_not), .in7(op3_not), .in8(op2_not), .in9(op1_not));
and10$ and_gate142(.out(and142), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8_not));
and10$ and_gate143(.out(and143), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not));
and9$ and_gate144(.out(and144), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op5_not), .in5(op4_not), .in6(op3_not), .in7(op2_not), .in8(op1));
and10$ and_gate145(.out(and145), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not));
and23$ and_gate146(.out(and146), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not), .in19(op5_not), .in20(op4_not), .in21(op3_not), .in22(op2_not));
and19$ and_gate147(.out(and147), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9), .in16(op8
), .in17(op7), .in18(op6));
and18$ and_gate148(.out(and148), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11), .in8(op10_not), .in9(op9_not), .in10(op8_not), .in11(op7_not), .in12(op6_not), .in13(op5_not), .in14(op4_not), .in15(op3_not), .in16(op2_not), .in17(op1_not));
and15$ and_gate149(.out(and149), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0), .in9(op10_not), .in10(op9), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not));
and16$ and_gate150(.out(and150), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4), .in13(op3), .in14(op2_not), .in15(op1_not));
and16$ and_gate151(.out(and151), .in0(sizeov_not), .in1(modrm7_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op8_not), .in9(op7), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and15$ and_gate152(.out(and152), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not));
and15$ and_gate153(.out(and153), .in0(modrm7_not), .in1(modrm6), .in2(modrm2_not), .in3(modrm1
), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13), .in8(op12_not), .in9(op8_not), .in10(op7_not), .in11(op6_not), .in12(op5_not), .in13(op4_not), .in14(op3));
and14$ and_gate154(.out(and154), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0), .in5(op15), .in6(op14), .in7(op13_not), .in8(op12_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and13$ and_gate155(.out(and155), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm0_not), .in4(op15), .in5(op14_not), .in6(op13
), .in7(op6_not), .in8(op5_not), .in9(op4_not), .in10(op3_not), .in11(op2_not), .in12(op1_not));
and13$ and_gate156(.out(and156), .in0(modrm3_not), .in1(modrm2), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not));
and10$ and_gate157(.out(and157), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not));
and9$ and_gate158(.out(and158), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9), .in8(op8));
and8$ and_gate159(.out(and159), .in0(sizeov), .in1(modrm7_not), .in2(modrm6
), .in3(op11), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op1_not));
and10$ and_gate160(.out(and160), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and9$ and_gate161(.out(and161), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op5_not), .in5(op4_not), .in6(op3_not), .in7(op2_not), .in8(op1));
and10$ and_gate162(.out(and162), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not));
and8$ and_gate163(.out(and163), .in0(op14), .in1(op13), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and8$ and_gate164(.out(and164), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1));
and23$ and_gate165(.out(and165), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not), .in19(op5_not), .in20(op4_not), .in21(op3_not), .in22(op2_not));
and17$ and_gate166(.out(and166), .in0(modrm1_not), .in1(modrm0_not), .in2(op15_not), .in3(op14_not), .in4(op13), .in5(op12), .in6(op11), .in7(op10
), .in8(op9), .in9(op8), .in10(op7), .in11(op6), .in12(op5), .in13(op4), .in14(op3_not), .in15(op2), .in16(op1_not));
and16$ and_gate167(.out(and167), .in0(sizeov), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(modrm4), .in5(modrm3), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1_not));
and16$ and_gate168(.out(and168), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8), .in9(op7), .in10(op6
), .in11(op5), .in12(op4), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and17$ and_gate169(.out(and169), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8));
and16$ and_gate170(.out(and170), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate171(.out(and171), .in0(sizeov), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate172(.out(and172), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and15$ and_gate173(.out(and173), .in0(modrm7_not), .in1(modrm6), .in2(modrm2_not), .in3(modrm1), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13), .in8(op12_not), .in9(op8_not), .in10(op7_not), .in11(op6_not), .in12(op5_not), .in13(op4_not), .in14(op3));
and15$ and_gate174(.out(and174), .in0(modrm6_not), .in1(modrm5), .in2(modrm1_not), .in3(modrm0), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not));
and13$ and_gate175(.out(and175), .in0(modrm3_not), .in1(modrm2), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13
), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not));
and14$ and_gate176(.out(and176), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and10$ and_gate177(.out(and177), .in0(modrm1_not), .in1(modrm0), .in2(op15), .in3(op14_not), .in4(op7), .in5(op6_not), .in6(op5), .in7(op4_not), .in8(op3), .in9(op2_not));
and10$ and_gate178(.out(and178), .in0(modrm3_not), .in1(modrm2), .in2(modrm1), .in3(modrm0_not), .in4(op9_not), .in5(op8_not), .in6(op7), .in7(op6_not), .in8(op5_not), .in9(op4_not));
and10$ and_gate179(.out(and179), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not));
and10$ and_gate180(.out(and180), .in0(modrm0), .in1(op15
), .in2(op14_not), .in3(op13_not), .in4(op6_not), .in5(op5_not), .in6(op4_not), .in7(op3_not), .in8(op2_not), .in9(op1_not));
and10$ and_gate181(.out(and181), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8_not));
and10$ and_gate182(.out(and182), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6
), .in3(modrm5), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and8$ and_gate183(.out(and183), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7));
and9$ and_gate184(.out(and184), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op5_not), .in5(op4_not), .in6(op3_not), .in7(op2_not), .in8(op1));
and10$ and_gate185(.out(and185), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not));
and8$ and_gate186(.out(and186), .in0(sizeov), .in1(op13), .in2(op12), .in3(op11_not), .in4(op10_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and8$ and_gate187(.out(and187), .in0(op14
), .in1(op13), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and8$ and_gate188(.out(and188), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1));
and23$ and_gate189(.out(and189), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5), .in4(modrm4), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6), .in19(op5_not), .in20(op4_not), .in21(op3_not), .in22(op1));
and21$ and_gate190(.out(and190), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(modrm1_not), .in5(modrm0
), .in6(op15_not), .in7(op14_not), .in8(op13_not), .in9(op12_not), .in10(op11_not), .in11(op10), .in12(op9_not), .in13(op8_not), .in14(op7), .in15(op6_not), .in16(op5_not), .in17(op4_not), .in18(op3_not), .in19(op2_not), .in20(op1_not));
and16$ and_gate191(.out(and191), .in0(modrm0_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7
), .in10(op6), .in11(op5), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not));
and18$ and_gate192(.out(and192), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8), .in17(op7));
and16$ and_gate193(.out(and193), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15), .in10(op14), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1));
and16$ and_gate194(.out(and194), .in0(
sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5), .in12(op4), .in13(op3), .in14(op2_not), .in15(op1_not));
and16$ and_gate195(.out(and195), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1), .in8(modrm0), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate196(.out(and196), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8
), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate197(.out(and197), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate198(.out(and198), .in0(sizeov_not), .in1(modrm7_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op8_not), .in9(op7), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate199(.out(and199), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and15$ and_gate200(.out(and200), .in0(modrm7_not), .in1(modrm6
), .in2(modrm2_not), .in3(modrm1), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13), .in8(op12_not), .in9(op8_not), .in10(op7_not), .in11(op6_not), .in12(op5_not), .in13(op4_not), .in14(op3));
and14$ and_gate201(.out(and201), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(modrm2_not), .in5(modrm1_not), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1));
and13$ and_gate202(.out(and202), .in0(modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(modrm1_not), .in5(modrm0), .in6(op7_not), .in7(op6_not), .in8(op5_not), .in9(op4_not), .in10(op3), .in11(op2), .in12(op1));
and14$ and_gate203(.out(and203), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10), .in10(op9), .in11(op8), .in12(op7_not), .in13(op6));
and15$ and_gate204(.out(and204), .in0(modrm6_not), .in1(modrm5), .in2(modrm1_not), .in3(modrm0), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not));
and14$ and_gate205(.out(and205), .in0(sizeov_not), .in1(op13_not), .in2(op12), .in3(op11), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7
), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate206(.out(and206), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0), .in5(op15), .in6(op14), .in7(op13_not), .in8(op12_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and13$ and_gate207(.out(and207), .in0(sizeov_not), .in1(modrm7), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op12), .in8(op11), .in9(op10_not), .in10(op9_not), .in11(op2_not), .in12(op1_not));
and13$ and_gate208(.out(and208), .in0(modrm3_not), .in1(modrm2), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not));
and10$ and_gate209(.out(and209), .in0(modrm2_not), .in1(modrm1), .in2(modrm0), .in3(op15_not), .in4(op8), .in5(op7_not), .in6(op6), .in7(op5_not), .in8(op4), .in9(op3_not));
and10$ and_gate210(.out(and210), .in0(modrm3_not), .in1(modrm2), .in2(modrm1), .in3(modrm0_not), .in4(op9_not), .in5(op8_not), .in6(op7), .in7(op6_not), .in8(op5_not), .in9(op4_not));
and10$ and_gate211(.out(and211), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and8$ and_gate212(.out(and212), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7));
and9$ and_gate213(.out(and213), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op5_not), .in5(op4_not), .in6(op3_not), .in7(op2_not), .in8(op1));
and8$ and_gate214(.out(and214), .in0(sizeov), .in1(op13), .in2(op12), .in3(op11_not), .in4(op10_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and24$ and_gate215(.out(and215), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3), .in6(modrm2_not), .in7(modrm1
), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not), .in19(op5_not), .in20(op4), .in21(op3), .in22(op2_not), .in23(op1_not));
and20$ and_gate216(.out(and216), .in0(modrm4_not), .in1(modrm3), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0_not), .in5(op15
), .in6(op14_not), .in7(op13_not), .in8(op12_not), .in9(op11_not), .in10(op10_not), .in11(op9), .in12(op8), .in13(op7_not), .in14(op6), .in15(op5), .in16(op4), .in17(op3), .in18(op2), .in19(op1));
and20$ and_gate217(.out(and217), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13_not), .in8(op12_not), .in9(op11_not), .in10(op10_not), .in11(op9), .in12(op8_not), .in13(op7_not), .in14(op6), .in15(op5_not), .in16(op4_not), .in17(op3_not), .in18(op2_not), .in19(op1_not));
and16$ and_gate218(.out(and218), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1));
and15$ and_gate219(.out(and219), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15_not), .in9(op14_not), .in10(op13), .in11(op7_not), .in12(op6), .in13(op2), .in14(op1));
and15$ and_gate220(.out(and220), .in0(modrm7), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5_not), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not));
and16$ and_gate221(.out(and221), .in0(sizeov
), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate222(.out(and222), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4), .in13(op3), .in14(op2_not), .in15(op1_not));
and16$ and_gate223(.out(and223), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate224(.out(and224), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and15$ and_gate225(.out(and225), .in0(modrm7_not), .in1(modrm6), .in2(modrm2_not), .in3(modrm1), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13), .in8(op12_not), .in9(op8_not), .in10(op7_not), .in11(op6_not), .in12(op5_not), .in13(op4_not), .in14(op3));
and14$ and_gate226(.out(and226), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(modrm2_not), .in5(modrm1_not), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1));
and14$ and_gate227(.out(and227), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10), .in10(op9), .in11(op8), .in12(op7_not), .in13(op6));
and15$ and_gate228(.out(and228), .in0(modrm6_not), .in1(modrm5), .in2(modrm1_not), .in3(modrm0), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not));
and14$ and_gate229(.out(and229), .in0(sizeov_not), .in1(op13_not), .in2(op12), .in3(op11), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate230(.out(and230), .in0(sizeov_not), .in1(modrm7_not), .in2(op12_not), .in3(op11), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and13$ and_gate231(.out(and231), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm0_not), .in4(op15), .in5(op14_not), .in6(op13
), .in7(op6_not), .in8(op5_not), .in9(op4_not), .in10(op3_not), .in11(op2_not), .in12(op1_not));
and13$ and_gate232(.out(and232), .in0(sizeov_not), .in1(modrm7), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op12), .in8(op11), .in9(op10_not), .in10(op9_not), .in11(op2_not), .in12(op1_not));
and10$ and_gate233(.out(and233), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5));
and10$ and_gate234(.out(and234), .in0(modrm1_not), .in1(modrm0
), .in2(op15), .in3(op14_not), .in4(op7), .in5(op6_not), .in6(op5), .in7(op4_not), .in8(op3), .in9(op2_not));
and8$ and_gate235(.out(and235), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(op11
), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op1_not));
and10$ and_gate236(.out(and236), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and8$ and_gate237(.out(and237), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(op10), .in5(op9
), .in6(op8_not), .in7(op7));
and10$ and_gate238(.out(and238), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not));
and21$ and_gate239(.out(and239), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(modrm1_not), .in5(modrm0), .in6(op15_not), .in7(op14_not), .in8(op13_not), .in9(op12_not), .in10(op11_not), .in11(op10), .in12(op9_not), .in13(op8_not), .in14(op7), .in15(op6_not), .in16(op5_not), .in17(op4_not), .in18(op3_not), .in19(op2_not), .in20(op1_not));
and19$ and_gate240(.out(and240), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9), .in16(op8), .in17(op7), .in18(op6));
and16$ and_gate241(.out(and241), .in0(sizeov), .in1(modrm7
), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4), .in13(op3_not), .in14(op2), .in15(op1_not));
and16$ and_gate242(.out(and242), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4), .in13(op3), .in14(op2_not), .in15(op1_not));
and14$ and_gate243(.out(and243), .in0(modrm6
), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(modrm2_not), .in5(modrm1_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3
), .in12(op2), .in13(op1));
and15$ and_gate244(.out(and244), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not));
and14$ and_gate245(.out(and245), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3), .in6(modrm2_not), .in7(modrm1), .in8(modrm0_not), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op1_not));
and15$ and_gate246(.out(and246), .in0(modrm7_not), .in1(modrm6), .in2(modrm2_not), .in3(modrm1), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13), .in8(op12_not), .in9(op8_not), .in10(op7_not), .in11(op6_not), .in12(op5_not), .in13(op4_not), .in14(op3));
and13$ and_gate247(.out(and247), .in0(modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(modrm1_not), .in5(modrm0
), .in6(op7_not), .in7(op6_not), .in8(op5_not), .in9(op4_not), .in10(op3), .in11(op2), .in12(op1));
and14$ and_gate248(.out(and248), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10), .in10(op9), .in11(op8), .in12(op7_not), .in13(op6));
and15$ and_gate249(.out(and249), .in0(modrm6_not), .in1(modrm5), .in2(modrm1_not), .in3(modrm0), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not));
and14$ and_gate250(.out(and250), .in0(sizeov_not), .in1(op13_not), .in2(op12), .in3(op11), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate251(.out(and251), .in0(sizeov_not), .in1(modrm7_not), .in2(op12_not), .in3(op11), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and13$ and_gate252(.out(and252), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm0_not), .in4(op15), .in5(op14_not), .in6(op13), .in7(op6_not), .in8(op5_not), .in9(op4_not), .in10(op3_not), .in11(op2_not), .in12(op1_not));
and14$ and_gate253(.out(and253), .in0(sizeov_not), .in1(modrm7
), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and13$ and_gate254(.out(and254), .in0(modrm3_not), .in1(modrm2), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not));
and11$ and_gate255(.out(and255), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4));
and10$ and_gate256(.out(and256), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5));
and8$ and_gate257(.out(and257), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(op11), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op1_not));
and8$ and_gate258(.out(and258), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7));
and9$ and_gate259(.out(and259), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op5_not), .in5(op4_not), .in6(op3_not), .in7(op2_not), .in8(op1));
and8$ and_gate260(.out(and260), .in0(sizeov), .in1(op13), .in2(op12), .in3(op11_not), .in4(op10_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and8$ and_gate261(.out(and261), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1));
and20$ and_gate262(.out(and262), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13_not), .in8(op12_not), .in9(op11_not), .in10(op10_not), .in11(op9), .in12(op8_not), .in13(op7_not), .in14(op6), .in15(op5_not), .in16(op4_not), .in17(op3_not), .in18(op2_not), .in19(op1_not));
and17$ and_gate263(.out(and263), .in0(
sizeov), .in1(modrm7), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8_not), .in12(op7), .in13(op6), .in14(op5), .in15(op4_not), .in16(op3));
and16$ and_gate264(.out(and264), .in0(sizeov_not), .in1(modrm7), .in2(modrm6
), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3), .in14(op2_not), .in15(op1));
and19$ and_gate265(.out(and265), .in0(modrm3_not), .in1(modrm2_not), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8), .in12(op7_not), .in13(op6_not), .in14(op5), .in15(op4_not), .in16(op3_not), .in17(op2_not), .in18(op1_not));
and15$ and_gate266(.out(and266), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not));
and14$ and_gate267(.out(and267), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10), .in10(op9), .in11(op8), .in12(op7_not), .in13(op6));
and15$ and_gate268(.out(and268), .in0(modrm6_not), .in1(modrm5), .in2(modrm1_not), .in3(modrm0), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not));
and14$ and_gate269(.out(and269), .in0(sizeov_not), .in1(modrm7_not), .in2(op12_not), .in3(op11), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate270(.out(and270), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(op9_not), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate271(.out(and271), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0
), .in5(op15), .in6(op14), .in7(op13_not), .in8(op12_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and11$ and_gate272(.out(and272), .in0(modrm3_not), .in1(modrm2
), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op5_not), .in7(op4), .in8(op3_not), .in9(op2), .in10(op1));
and13$ and_gate273(.out(and273), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm0_not), .in4(op15), .in5(op14_not), .in6(op13), .in7(op6_not), .in8(op5_not), .in9(op4_not), .in10(op3_not), .in11(op2_not), .in12(op1_not));
and13$ and_gate274(.out(and274), .in0(sizeov_not), .in1(modrm7), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op12), .in8(op11), .in9(op10_not), .in10(op9_not), .in11(op2_not), .in12(op1_not));
and11$ and_gate275(.out(and275), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2
), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4));
and10$ and_gate276(.out(and276), .in0(modrm2_not), .in1(modrm1), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13), .in6(op4_not), .in7(op3), .in8(op2), .in9(op1_not));
and10$ and_gate277(.out(and277), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3), .in6(op8
), .in7(op7), .in8(op6_not), .in9(op5));
and10$ and_gate278(.out(and278), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13), .in6(op4_not), .in7(op3_not), .in8(op2), .in9(op1_not));
and8$ and_gate279(.out(and279), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7));
and10$ and_gate280(.out(and280), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not));
and8$ and_gate281(.out(and281), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1));
and17$ and_gate282(.out(and282), .in0(sizeov), .in1(modrm7), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1
), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8_not), .in12(op7), .in13(op6), .in14(op5), .in15(op4_not), .in16(op3));
and19$ and_gate283(.out(and283), .in0(modrm3_not), .in1(modrm2_not), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8), .in12(op7_not), .in13(op6_not), .in14(op5), .in15(op4_not), .in16(op3_not), .in17(op2_not), .in18(op1_not));
and16$ and_gate284(.out(and284), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5
), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15), .in10(op14), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1));
and16$ and_gate285(.out(and285), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4), .in13(op3), .in14(op2_not), .in15(op1_not));
and16$ and_gate286(.out(and286), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and13$ and_gate287(.out(and287), .in0(sizeov_not), .in1(modrm7), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2), .in7(modrm1_not), .in8(modrm0
), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2));
and13$ and_gate288(.out(and288), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0), .in5(op15_not), .in6(op14_not), .in7(op13), .in8(op12), .in9(op11_not), .in10(op10), .in11(op9_not), .in12(op8));
and15$ and_gate289(.out(and289), .in0(modrm7_not), .in1(modrm6), .in2(modrm2_not), .in3(modrm1), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13), .in8(op12_not), .in9(op8_not), .in10(op7_not), .in11(op6_not), .in12(op5_not), .in13(op4_not), .in14(op3));
and14$ and_gate290(.out(and290), .in0(
sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate291(.out(and291), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(modrm2_not), .in5(modrm1_not), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1));
and14$ and_gate292(.out(and292), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10), .in10(op9), .in11(op8), .in12(op7_not), .in13(op6));
and14$ and_gate293(.out(and293), .in0(sizeov_not), .in1(op13_not), .in2(op12), .in3(op11), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate294(.out(and294), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(op9_not), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and11$ and_gate295(.out(and295), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4
), .in5(modrm3_not), .in6(modrm2), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4));
and10$ and_gate296(.out(and296), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5
), .in4(modrm4_not), .in5(modrm3), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5));
and8$ and_gate297(.out(and297), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1));
and20$ and_gate298(.out(and298), .in0(modrm4_not), .in1(modrm3), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0_not), .in5(op15), .in6(op14_not), .in7(op13_not), .in8(op12_not), .in9(op11_not), .in10(op10_not), .in11(op9), .in12(op8), .in13(op7_not), .in14(op6), .in15(op5), .in16(op4), .in17(op3), .in18(op2), .in19(op1));
and21$ and_gate299(.out(and299), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(modrm1_not), .in5(modrm0), .in6(op15_not), .in7(op14_not), .in8(op13_not), .in9(op12_not), .in10(op11_not), .in11(op10
), .in12(op9_not), .in13(op8_not), .in14(op7), .in15(op6_not), .in16(op5_not), .in17(op4_not), .in18(op3_not), .in19(op2_not), .in20(op1_not));
and20$ and_gate300(.out(and300), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0), .in5(op15_not), .in6(op14_not), .in7(op13), .in8(op12_not), .in9(op11_not), .in10(op10_not), .in11(op9_not), .in12(op8_not), .in13(op7_not), .in14(op6_not), .in15(op5_not), .in16(op4_not), .in17(op3_not), .in18(op2_not), .in19(op1_not));
and17$ and_gate301(.out(and301), .in0(sizeov), .in1(modrm7), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8_not), .in12(op7), .in13(op6), .in14(op5), .in15(op4_not), .in16(op3));
and16$ and_gate302(.out(and302), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and15$ and_gate303(.out(and303), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not));
and13$ and_gate304(.out(and304), .in0(sizeov_not), .in1(modrm7), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2), .in7(modrm1_not), .in8(modrm0
), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2));
and15$ and_gate305(.out(and305), .in0(modrm7_not), .in1(modrm6), .in2(modrm2_not), .in3(modrm1), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13), .in8(op12_not), .in9(op8_not), .in10(op7_not), .in11(op6_not), .in12(op5_not), .in13(op4_not), .in14(op3));
and14$ and_gate306(.out(and306), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and15$ and_gate307(.out(and307), .in0(modrm6_not), .in1(modrm5), .in2(modrm1_not), .in3(modrm0), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not));
and14$ and_gate308(.out(and308), .in0(sizeov_not), .in1(op13_not), .in2(op12), .in3(op11), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7
), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate309(.out(and309), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op11_not), .in4(op10
), .in5(op9), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not));
and14$ and_gate310(.out(and310), .in0(sizeov_not), .in1(modrm7_not), .in2(op12_not), .in3(op11), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate311(.out(and311), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(op9_not), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate312(.out(and312), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and11$ and_gate313(.out(and313), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4));
and10$ and_gate314(.out(and314), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5));
and10$ and_gate315(.out(and315), .in0(sizeov), .in1(modrm7_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11), .in8(op2_not), .in9(op1_not));
and10$ and_gate316(.out(and316), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13), .in6(op4_not), .in7(op3_not), .in8(op2), .in9(op1_not));
and10$ and_gate317(.out(and317), .in0(sizeov_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op3_not), .in8(op2_not), .in9(op1));
and8$ and_gate318(.out(and318), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5
), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7));
and8$ and_gate319(.out(and319), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1));
and20$ and_gate320(.out(and320), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13_not), .in8(op12_not), .in9(op11_not), .in10(op10_not), .in11(op9), .in12(op8_not), .in13(op7_not), .in14(op6), .in15(op5_not), .in16(op4_not), .in17(op3_not), .in18(op2_not), .in19(op1_not));
and19$ and_gate321(.out(and321), .in0(modrm3_not), .in1(modrm2_not), .in2(modrm1_not), .in3(modrm0_not), .in4(op15), .in5(op14_not), .in6(op13), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8_not), .in12(op7_not), .in13(op6_not), .in14(op5_not), .in15(op4_not), .in16(op3_not), .in17(op2_not), .in18(op1_not));
and17$ and_gate322(.out(and322), .in0(sizeov), .in1(modrm7), .in2(modrm6
), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8_not), .in12(op7), .in13(op6
), .in14(op5), .in15(op4_not), .in16(op3));
and13$ and_gate323(.out(and323), .in0(sizeov_not), .in1(modrm7), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2
), .in7(modrm1_not), .in8(modrm0), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2));
and14$ and_gate324(.out(and324), .in0(sizeov), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate325(.out(and325), .in0(
sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate326(.out(and326), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(modrm2_not), .in5(modrm1_not), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1));
and14$ and_gate327(.out(and327), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10), .in10(op9), .in11(op8), .in12(op7_not), .in13(op6));
and15$ and_gate328(.out(and328), .in0(modrm6_not), .in1(modrm5), .in2(modrm1_not), .in3(modrm0), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not));
and14$ and_gate329(.out(and329), .in0(sizeov_not), .in1(op13_not), .in2(op12), .in3(op11), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7
), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate330(.out(and330), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op10_not), .in5(op9), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate331(.out(and331), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op11_not), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not));
and13$ and_gate332(.out(and332), .in0(sizeov_not), .in1(modrm7), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op12), .in8(op11), .in9(op10_not), .in10(op9_not), .in11(op2_not), .in12(op1_not));
and14$ and_gate333(.out(and333), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and11$ and_gate334(.out(and334), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4));
and11$ and_gate335(.out(and335), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14), .in5(op13), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op9_not), .in10(op8));
and9$ and_gate336(.out(and336), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9), .in8(op8));
and10$ and_gate337(.out(and337), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op1_not));
and8$ and_gate338(.out(and338), .in0(sizeov), .in1(op13), .in2(op12), .in3(op11_not), .in4(op10_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and21$ and_gate339(.out(and339), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(modrm1_not), .in5(modrm0), .in6(op15_not), .in7(op14_not), .in8(op13_not), .in9(op12_not), .in10(op11_not), .in11(op10), .in12(op9_not), .in13(op8_not), .in14(op7), .in15(op6_not), .in16(op5_not), .in17(op4_not), .in18(op3_not), .in19(op2_not), .in20(op1_not));
and17$ and_gate340(.out(and340), .in0(
sizeov), .in1(modrm7), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8_not), .in12(op7), .in13(op6), .in14(op5), .in15(op4_not), .in16(op3));
and18$ and_gate341(.out(and341), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8), .in17(op7));
and18$ and_gate342(.out(and342), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11), .in8(op10_not), .in9(op9_not), .in10(op8_not), .in11(op7_not), .in12(op6_not), .in13(op5_not), .in14(op4_not), .in15(op3_not), .in16(op2_not), .in17(op1_not));
and15$ and_gate343(.out(and343), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0), .in9(op10_not), .in10(op9), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not));
and13$ and_gate344(.out(and344), .in0(sizeov_not), .in1(modrm7
), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2), .in7(modrm1_not), .in8(modrm0), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2));
and14$ and_gate345(.out(and345), .in0(
sizeov), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate346(.out(and346), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op10_not), .in5(op9
), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate347(.out(and347), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op11_not), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not));
and14$ and_gate348(.out(and348), .in0(sizeov_not), .in1(modrm7_not), .in2(op12_not), .in3(op11), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate349(.out(and349), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(op9_not), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and13$ and_gate350(.out(and350), .in0(sizeov_not), .in1(modrm7), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13
), .in7(op12), .in8(op11), .in9(op10_not), .in10(op9_not), .in11(op2_not), .in12(op1_not));
and14$ and_gate351(.out(and351), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and13$ and_gate352(.out(and352), .in0(modrm3_not), .in1(modrm2), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not));
and10$ and_gate353(.out(and353), .in0(sizeov_not), .in1(modrm1_not), .in2(modrm0), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op3_not), .in8(op2), .in9(op1));
and9$ and_gate354(.out(and354), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9), .in8(op8));
and10$ and_gate355(.out(and355), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and17$ and_gate356(.out(and356), .in0(modrm1_not), .in1(modrm0_not), .in2(op15_not), .in3(op14_not), .in4(op13), .in5(op12), .in6(op11), .in7(op10), .in8(op9), .in9(op8), .in10(op7
), .in11(op6), .in12(op5), .in13(op4), .in14(op3_not), .in15(op2), .in16(op1_not));
and20$ and_gate357(.out(and357), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13_not), .in8(op12_not), .in9(op11_not), .in10(op10_not), .in11(op9), .in12(op8_not), .in13(op7_not), .in14(op6), .in15(op5_not), .in16(op4_not), .in17(op3_not), .in18(op2_not), .in19(op1_not));
and16$ and_gate358(.out(and358), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5), .in12(op4), .in13(op3), .in14(op2_not), .in15(op1_not));
and16$ and_gate359(.out(and359), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6
), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15), .in10(op9_not), .in11(op8), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and15$ and_gate360(.out(and360), .in0(modrm7), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6), .in10(op5_not), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not));
and16$ and_gate361(.out(and361), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6
), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and13$ and_gate362(.out(and362), .in0(sizeov_not), .in1(modrm7), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2), .in7(modrm1_not), .in8(modrm0
), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2));
and14$ and_gate363(.out(and363), .in0(sizeov), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate364(.out(and364), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate365(.out(and365), .in0(
sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op10_not), .in5(op9), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate366(.out(and366), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op11_not), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7_not), .in8(op6
), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not));
and14$ and_gate367(.out(and367), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and11$ and_gate368(.out(and368), .in0(sizeov_not), .in1(modrm7
), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4));
and14$ and_gate369(.out(and369), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and10$ and_gate370(.out(and370), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm0_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op2_not), .in9(op1_not));
and10$ and_gate371(.out(and371), .in0(sizeov_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op3_not), .in8(op2_not), .in9(op1));
and10$ and_gate372(.out(and372), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and8$ and_gate373(.out(and373), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(op11), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op1_not));
and10$ and_gate374(.out(and374), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not));
and21$ and_gate375(.out(and375), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1
), .in8(modrm0_not), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8), .in17(op7_not), .in18(op3), .in19(op2), .in20(op1));
and23$ and_gate376(.out(and376), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not), .in19(op5_not), .in20(op4_not), .in21(op3_not), .in22(op2_not));
and22$ and_gate377(.out(and377), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not), .in19(op5_not), .in20(op4_not), .in21(op3_not));
and17$ and_gate378(.out(and378), .in0(sizeov), .in1(modrm7), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8_not), .in12(op7), .in13(op6), .in14(op5), .in15(op4_not), .in16(op3));
and16$ and_gate379(.out(and379), .in0(modrm0_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4), .in13(op3
), .in14(op2), .in15(op1_not));
and19$ and_gate380(.out(and380), .in0(modrm3_not), .in1(modrm2_not), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8), .in12(op7_not), .in13(op6_not), .in14(op5), .in15(op4_not), .in16(op3_not), .in17(op2_not), .in18(op1_not));
and16$ and_gate381(.out(and381), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1), .in8(modrm0), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and14$ and_gate382(.out(and382), .in0(modrm6), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(modrm2_not), .in5(modrm1_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3), .in12(op2), .in13(op1));
and14$ and_gate383(.out(and383), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10), .in10(op9), .in11(op8
), .in12(op7_not), .in13(op6));
and14$ and_gate384(.out(and384), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op10_not), .in5(op9), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate385(.out(and385), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op11_not), .in4(op10), .in5(op9
), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not));
and14$ and_gate386(.out(and386), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(op9_not), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate387(.out(and387), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(op7_not), .in8(op6), .in9(op5
), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate388(.out(and388), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and10$ and_gate389(.out(and389), .in0(
sizeov), .in1(modrm7_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11), .in8(op2_not), .in9(op1_not));
and10$ and_gate390(.out(and390), .in0(sizeov_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op3_not), .in8(op2_not), .in9(op1));
and10$ and_gate391(.out(and391), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op15_not), .in4(op14), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op1_not));
and20$ and_gate392(.out(and392), .in0(modrm4_not), .in1(modrm3), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0_not), .in5(op15), .in6(op14_not), .in7(op13_not), .in8(op12_not), .in9(op11_not), .in10(op10_not), .in11(op9), .in12(op8), .in13(op7_not), .in14(op6), .in15(op5), .in16(op4), .in17(op3), .in18(op2), .in19(op1));
and22$ and_gate393(.out(and393), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not), .in19(op5_not), .in20(op4_not), .in21(op3_not));
and17$ and_gate394(.out(and394), .in0(modrm1_not), .in1(modrm0_not), .in2(op15_not), .in3(op14_not), .in4(op13), .in5(op12), .in6(op11), .in7(op10), .in8(op9), .in9(op8), .in10(op7), .in11(op6), .in12(op5
), .in13(op4), .in14(op3_not), .in15(op2), .in16(op1_not));
and16$ and_gate395(.out(and395), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9
), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1));
and18$ and_gate396(.out(and396), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11), .in8(op10_not), .in9(op9_not), .in10(op8_not), .in11(op7_not), .in12(op6_not), .in13(op5_not), .in14(op4_not), .in15(op3_not), .in16(op2_not), .in17(op1_not));
and16$ and_gate397(.out(and397), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0), .in9(op15), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11), .in14(op2_not), .in15(op1_not));
and15$ and_gate398(.out(and398), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15_not), .in9(op14_not), .in10(op13), .in11(op7_not), .in12(op6), .in13(op2), .in14(op1));
and14$ and_gate399(.out(and399), .in0(sizeov), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and15$ and_gate400(.out(and400), .in0(modrm6_not), .in1(modrm5), .in2(modrm1_not), .in3(modrm0), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not));
and14$ and_gate401(.out(and401), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op10_not), .in5(op9), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate402(.out(and402), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(op9_not), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate403(.out(and403), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate404(.out(and404), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and10$ and_gate405(.out(and405), .in0(sizeov), .in1(modrm7_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11), .in8(op2_not), .in9(op1_not));
and10$ and_gate406(.out(and406), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13), .in6(op4_not), .in7(op3_not), .in8(op2), .in9(op1_not));
and10$ and_gate407(.out(and407), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op14_not), .in5(op13), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate408(.out(and408), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op1_not));
and10$ and_gate409(.out(and409), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate410(.out(and410), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not));
and16$ and_gate411(.out(and411), .in0(modrm0_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5
), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not));
and16$ and_gate412(.out(and412), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3
), .in6(modrm2_not), .in7(modrm1), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12), .in13(op6_not), .in14(op5), .in15(op1));
and15$ and_gate413(.out(and413), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0
), .in9(op10_not), .in10(op9), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not));
and14$ and_gate414(.out(and414), .in0(modrm6), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(modrm2_not), .in5(modrm1_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3), .in12(op2), .in13(op1));
and14$ and_gate415(.out(and415), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3), .in6(modrm2_not), .in7(modrm1), .in8(modrm0_not), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op1_not));
and14$ and_gate416(.out(and416), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate417(.out(and417), .in0(sizeov_not), .in1(modrm7
), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate418(.out(and418), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and10$ and_gate419(.out(and419), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op1_not));
and10$ and_gate420(.out(and420), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8_not));
and10$ and_gate421(.out(and421), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not));
and10$ and_gate422(.out(and422), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not));
and21$ and_gate423(.out(and423), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1
), .in8(modrm0_not), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8), .in17(op7_not), .in18(op3), .in19(op2), .in20(op1));
and23$ and_gate424(.out(and424), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not), .in19(op5_not), .in20(op4_not), .in21(op3_not), .in22(op2_not));
and17$ and_gate425(.out(and425), .in0(sizeov), .in1(modrm7), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8_not), .in12(op7), .in13(op6), .in14(op5), .in15(op4_not), .in16(op3));
and16$ and_gate426(.out(and426), .in0(modrm0_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not));
and16$ and_gate427(.out(and427), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1));
and16$ and_gate428(.out(and428), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14), .in11(op13), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9));
and16$ and_gate429(.out(and429), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15), .in10(op9_not), .in11(op8), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and14$ and_gate430(.out(and430), .in0(sizeov), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate431(.out(and431), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(op7_not), .in8(op6), .in9(op5
), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and11$ and_gate432(.out(and432), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4));
and14$ and_gate433(.out(and433), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and10$ and_gate434(.out(and434), .in0(modrm3_not), .in1(modrm2), .in2(modrm1), .in3(modrm0_not), .in4(op9_not), .in5(op8_not), .in6(op7), .in7(op6_not), .in8(op5_not), .in9(op4_not));
and21$ and_gate435(.out(and435), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1
), .in8(modrm0_not), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8), .in17(op7_not), .in18(op3), .in19(op2), .in20(op1));
and17$ and_gate436(.out(and436), .in0(
sizeov), .in1(modrm7), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8_not), .in12(op7), .in13(op6), .in14(op5), .in15(op4_not), .in16(op3));
and16$ and_gate437(.out(and437), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1));
and17$ and_gate438(.out(and438), .in0(sizeov
), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15
), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8));
and16$ and_gate439(.out(and439), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1), .in8(modrm0), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12
), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate440(.out(and440), .in0(sizeov), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and15$ and_gate441(.out(and441), .in0(modrm7_not), .in1(modrm6), .in2(modrm2_not), .in3(modrm1), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13), .in8(op12_not), .in9(op8_not), .in10(op7_not), .in11(op6_not), .in12(op5_not), .in13(op4_not), .in14(op3));
and13$ and_gate442(.out(and442), .in0(modrm3_not), .in1(modrm2), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not));
and14$ and_gate443(.out(and443), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and10$ and_gate444(.out(and444), .in0(modrm2_not), .in1(modrm1), .in2(modrm0
), .in3(op15_not), .in4(op8), .in5(op7_not), .in6(op6), .in7(op5_not), .in8(op4), .in9(op3_not));
and10$ and_gate445(.out(and445), .in0(sizeov_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op3_not), .in8(op2_not), .in9(op1));
and10$ and_gate446(.out(and446), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not));
and16$ and_gate447(.out(and447), .in0(sizeov), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(modrm4), .in5(modrm3), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1_not));
and18$ and_gate448(.out(and448), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9), .in16(op3_not), .in17(op2));
and18$ and_gate449(.out(and449), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8), .in17(op7));
and16$ and_gate450(.out(and450), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0), .in9(op15), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11), .in14(op2_not), .in15(op1_not));
and16$ and_gate451(.out(and451), .in0(sizeov_not), .in1(modrm7_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op8_not), .in9(op7), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and13$ and_gate452(.out(and452), .in0(sizeov_not), .in1(modrm7), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2), .in7(modrm1_not), .in8(modrm0), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2));
and14$ and_gate453(.out(and453), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op11_not), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not));
and13$ and_gate454(.out(and454), .in0(modrm3_not), .in1(modrm2), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not));
and10$ and_gate455(.out(and455), .in0(
sizeov), .in1(modrm7_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11), .in8(op2_not), .in9(op1_not));
and10$ and_gate456(.out(and456), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not));
and19$ and_gate457(.out(and457), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not));
and16$ and_gate458(.out(and458), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15), .in10(op9_not), .in11(op8), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate459(.out(and459), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1), .in8(modrm0), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and15$ and_gate460(.out(and460), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15_not), .in9(op14_not), .in10(op13), .in11(op7_not), .in12(op6), .in13(op2), .in14(op1));
and16$ and_gate461(.out(and461), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6
), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and14$ and_gate462(.out(and462), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3), .in6(modrm2_not), .in7(modrm1), .in8(modrm0_not), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op1_not));
and15$ and_gate463(.out(and463), .in0(modrm7_not), .in1(modrm6), .in2(modrm2_not), .in3(modrm1), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13), .in8(op12_not), .in9(op8_not), .in10(op7_not), .in11(op6_not), .in12(op5_not), .in13(op4_not), .in14(op3));
and14$ and_gate464(.out(and464), .in0(sizeov
), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op10_not), .in5(op9), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate465(.out(and465), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op11_not), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5
), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not));
and14$ and_gate466(.out(and466), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and11$ and_gate467(.out(and467), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14), .in5(op13), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op9_not), .in10(op8));
and10$ and_gate468(.out(and468), .in0(modrm1_not), .in1(modrm0), .in2(op15), .in3(op14_not), .in4(op7), .in5(op6_not), .in6(op5), .in7(op4_not), .in8(op3), .in9(op2_not));
and10$ and_gate469(.out(and469), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op1_not));
and10$ and_gate470(.out(and470), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not));
and24$ and_gate471(.out(and471), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3), .in6(modrm2_not), .in7(modrm1
), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not), .in19(op5_not), .in20(op4), .in21(op3), .in22(op2_not), .in23(op1_not));
and18$ and_gate472(.out(and472), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9), .in16(op3_not), .in17(op2));
and19$ and_gate473(.out(and473), .in0(modrm3_not), .in1(modrm2_not), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8), .in12(op7_not), .in13(op6_not), .in14(op5), .in15(op4_not), .in16(op3_not), .in17(op2_not), .in18(op1_not));
and16$ and_gate474(.out(and474), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14
), .in11(op13), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9));
and16$ and_gate475(.out(and475), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3), .in6(modrm2_not), .in7(modrm1), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12), .in13(op6_not), .in14(op5), .in15(op1));
and16$ and_gate476(.out(and476), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0), .in9(op15), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11), .in14(op2_not), .in15(op1_not));
and15$ and_gate477(.out(and477), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3), .in5(modrm2), .in6(modrm1_not), .in7(modrm0_not), .in8(op15_not), .in9(op14_not), .in10(op13), .in11(op7_not), .in12(op6), .in13(op2), .in14(op1));
and16$ and_gate478(.out(and478), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and14$ and_gate479(.out(and479), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3), .in6(modrm2_not), .in7(modrm1), .in8(modrm0_not), .in9(op15_not), .in10(op14
), .in11(op13_not), .in12(op12_not), .in13(op1_not));
and14$ and_gate480(.out(and480), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op11_not), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not));
and11$ and_gate481(.out(and481), .in0(modrm1_not), .in1(modrm0_not), .in2(op15_not), .in3(op14), .in4(op13_not), .in5(op12
), .in6(op11_not), .in7(op10_not), .in8(op9), .in9(op8_not), .in10(op7));
and11$ and_gate482(.out(and482), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14), .in5(op13
), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op9_not), .in10(op8));
and10$ and_gate483(.out(and483), .in0(sizeov_not), .in1(modrm1_not), .in2(modrm0), .in3(op15_not), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op3_not), .in8(op2), .in9(op1));
and10$ and_gate484(.out(and484), .in0(modrm1_not), .in1(modrm0), .in2(op15), .in3(op14_not), .in4(op7), .in5(op6_not), .in6(op5
), .in7(op4_not), .in8(op3), .in9(op2_not));
and10$ and_gate485(.out(and485), .in0(modrm0), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op6_not), .in5(op5_not), .in6(op4_not), .in7(op3_not), .in8(op2_not), .in9(op1_not));
and10$ and_gate486(.out(and486), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not));
and10$ and_gate487(.out(and487), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not));
and9$ and_gate488(.out(and488), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op5_not), .in5(op4_not), .in6(op3_not), .in7(op2_not), .in8(op1));
and18$ and_gate489(.out(and489), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9), .in16(op3_not), .in17(op2));
and16$ and_gate490(.out(and490), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3), .in6(modrm2_not), .in7(modrm1), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12), .in13(op6_not), .in14(op5), .in15(op1));
and16$ and_gate491(.out(and491), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0), .in9(op15), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11
), .in14(op2_not), .in15(op1_not));
and16$ and_gate492(.out(and492), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4), .in13(op3), .in14(op2_not), .in15(op1_not));
and16$ and_gate493(.out(and493), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and13$ and_gate494(.out(and494), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0), .in5(op15_not), .in6(op14_not), .in7(op13), .in8(op12), .in9(op11_not), .in10(op10), .in11(op9_not), .in12(op8));
and14$ and_gate495(.out(and495), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op10_not), .in5(op9), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate496(.out(and496), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0), .in5(op15), .in6(op14), .in7(op13_not), .in8(op12_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and11$ and_gate497(.out(and497), .in0(modrm1_not), .in1(modrm0_not), .in2(op15_not), .in3(op14), .in4(op13_not), .in5(op12), .in6(op11_not), .in7(op10_not), .in8(op9), .in9(op8_not), .in10(op7));
and10$ and_gate498(.out(and498), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13), .in6(op4_not), .in7(op3_not), .in8(op2), .in9(op1_not));
and10$ and_gate499(.out(and499), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op14_not), .in5(op13), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate500(.out(and500), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op15_not), .in4(op14), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op1_not));
and10$ and_gate501(.out(and501), .in0(
modrm0), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op6_not), .in5(op5_not), .in6(op4_not), .in7(op3_not), .in8(op2_not), .in9(op1_not));
and9$ and_gate502(.out(and502), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op5_not), .in5(op4_not), .in6(op3_not), .in7(op2_not), .in8(op1));
and8$ and_gate503(.out(and503), .in0(op14), .in1(op13), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and18$ and_gate504(.out(and504), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0), .in9(op15_not), .in10(op14), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9), .in16(op3_not), .in17(op2));
and16$ and_gate505(.out(and505), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3), .in6(modrm2_not), .in7(modrm1), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12), .in13(op6_not), .in14(op5), .in15(op1));
and15$ and_gate506(.out(and506), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(modrm3_not), .in5(modrm2), .in6(op9_not), .in7(op8_not), .in8(op7), .in9(op6_not), .in10(op5_not), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not));
and15$ and_gate507(.out(and507), .in0(modrm6_not), .in1(modrm5), .in2(modrm1_not), .in3(modrm0), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not));
and14$ and_gate508(.out(and508), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0), .in5(op15
), .in6(op14), .in7(op13_not), .in8(op12_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and10$ and_gate509(.out(and509), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op15_not), .in4(op14), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op1_not));
and10$ and_gate510(.out(and510), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9_not), .in8(op8_not), .in9(op7_not));
and10$ and_gate511(.out(and511), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8_not));
and8$ and_gate512(.out(and512), .in0(sizeov), .in1(op13), .in2(op12), .in3(op11_not), .in4(op10_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and8$ and_gate513(.out(and513), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1));
and21$ and_gate514(.out(and514), .in0(sizeov), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(modrm4), .in5(modrm3), .in6(modrm2), .in7(modrm1
), .in8(modrm0), .in9(op15), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10), .in15(op9), .in16(op8), .in17(op7_not), .in18(op6), .in19(op5), .in20(op4_not));
and23$ and_gate515(.out(and515), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not), .in19(op5_not), .in20(op4_not), .in21(op3_not), .in22(op2_not));
and14$ and_gate516(.out(and516), .in0(modrm6_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(modrm2_not), .in5(modrm1_not), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3), .in12(op2_not), .in13(op1));
and14$ and_gate517(.out(and517), .in0(sizeov_not), .in1(op13_not), .in2(op12), .in3(op11), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate518(.out(and518), .in0(sizeov_not), .in1(modrm7_not), .in2(op12_not), .in3(op11), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and13$ and_gate519(.out(and519), .in0(sizeov_not), .in1(modrm7), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op12), .in8(op11), .in9(op10_not), .in10(op9_not), .in11(op2_not), .in12(op1_not));
and13$ and_gate520(.out(and520), .in0(modrm3_not), .in1(modrm2), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not));
and10$ and_gate521(.out(and521), .in0(modrm1_not), .in1(modrm0), .in2(op15), .in3(op14_not), .in4(op7), .in5(op6_not), .in6(op5), .in7(op4_not), .in8(op3), .in9(op2_not));
and8$ and_gate522(.out(and522), .in0(sizeov), .in1(op13), .in2(op12), .in3(op11_not), .in4(op10_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and8$ and_gate523(.out(and523), .in0(op14
), .in1(op13), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and8$ and_gate524(.out(and524), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1));
and22$ and_gate525(.out(and525), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not), .in19(op5_not), .in20(op4_not), .in21(op3_not));
and21$ and_gate526(.out(and526), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(modrm2_not), .in4(modrm1_not), .in5(modrm0), .in6(op15_not), .in7(op14_not), .in8(op13_not), .in9(op12_not), .in10(op11_not), .in11(op10), .in12(op9_not), .in13(op8_not), .in14(op7), .in15(op6_not), .in16(op5_not), .in17(op4_not), .in18(op3_not), .in19(op2_not), .in20(op1_not));
and16$ and_gate527(.out(and527), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and15$ and_gate528(.out(and528), .in0(modrm7_not), .in1(modrm6
), .in2(modrm2_not), .in3(modrm1), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13), .in8(op12_not), .in9(op8_not), .in10(op7_not), .in11(op6_not), .in12(op5_not), .in13(op4_not), .in14(op3));
and14$ and_gate529(.out(and529), .in0(sizeov_not), .in1(op13_not), .in2(op12), .in3(op11), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate530(.out(and530), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op11_not), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not));
and13$ and_gate531(.out(and531), .in0(sizeov_not), .in1(modrm7), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op12), .in8(op11), .in9(op10_not), .in10(op9_not), .in11(op2_not), .in12(op1_not));
and11$ and_gate532(.out(and532), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14), .in5(op13), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op9_not), .in10(op8));
and10$ and_gate533(.out(and533), .in0(modrm7_not), .in1(modrm6_not), .in2(modrm5_not), .in3(modrm4_not), .in4(op13_not), .in5(op12), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8_not));
and10$ and_gate534(.out(and534), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(op10_not), .in5(op9_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not));
and8$ and_gate535(.out(and535), .in0(sizeov), .in1(op13), .in2(op12
), .in3(op11_not), .in4(op10_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and21$ and_gate536(.out(and536), .in0(sizeov), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(modrm4), .in5(modrm3), .in6(modrm2), .in7(modrm1
), .in8(modrm0), .in9(op15), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10), .in15(op9), .in16(op8), .in17(op7_not), .in18(op6), .in19(op5), .in20(op4_not));
and20$ and_gate537(.out(and537), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0_not), .in5(op15_not), .in6(op14_not), .in7(op13_not), .in8(op12_not), .in9(op11_not), .in10(op10_not), .in11(op9), .in12(op8_not), .in13(op7_not), .in14(op6), .in15(op5_not), .in16(op4_not), .in17(op3_not), .in18(op2_not), .in19(op1_not));
and16$ and_gate538(.out(and538), .in0(sizeov_not), .in1(modrm7
), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4), .in13(op3_not), .in14(op2), .in15(op1_not));
and13$ and_gate539(.out(and539), .in0(modrm0_not), .in1(op15_not), .in2(op14), .in3(op13_not), .in4(op12), .in5(op11_not), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4));
and14$ and_gate540(.out(and540), .in0(
sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op10_not), .in5(op9), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate541(.out(and541), .in0(sizeov_not), .in1(modrm7_not), .in2(op12_not), .in3(op11), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate542(.out(and542), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0), .in5(op15
), .in6(op14), .in7(op13_not), .in8(op12_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and13$ and_gate543(.out(and543), .in0(sizeov_not), .in1(modrm7), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13), .in7(op12), .in8(op11), .in9(op10_not), .in10(op9_not), .in11(op2_not), .in12(op1_not));
and11$ and_gate544(.out(and544), .in0(modrm1_not), .in1(modrm0_not), .in2(op15_not), .in3(op14), .in4(op13_not), .in5(op12), .in6(op11_not), .in7(op10_not), .in8(op9), .in9(op8_not), .in10(op7));
and11$ and_gate545(.out(and545), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14), .in5(op13), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op9_not), .in10(op8));
and10$ and_gate546(.out(and546), .in0(modrm1_not), .in1(modrm0), .in2(op15), .in3(op14_not), .in4(op7), .in5(op6_not), .in6(op5), .in7(op4_not), .in8(op3), .in9(op2_not));
and8$ and_gate547(.out(and547), .in0(sizeov
), .in1(modrm7_not), .in2(modrm6), .in3(op11), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op1_not));
and8$ and_gate548(.out(and548), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1));
and20$ and_gate549(.out(and549), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3), .in6(modrm2
), .in7(modrm1), .in8(modrm0), .in9(op15_not), .in10(op14_not), .in11(op13), .in12(op12_not), .in13(op11), .in14(op10), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6
), .in19(op5));
and22$ and_gate550(.out(and550), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13_not), .in12(op12_not), .in13(op11_not), .in14(op10), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6_not), .in19(op5_not), .in20(op4_not), .in21(op3_not));
and19$ and_gate551(.out(and551), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2_not), .in7(modrm1_not), .in8(modrm0_not), .in9(op15_not), .in10(op14_not), .in11(op13), .in12(op12_not), .in13(op11_not), .in14(op10_not), .in15(op9), .in16(op8), .in17(op7), .in18(op6));
and19$ and_gate552(.out(and552), .in0(modrm3_not), .in1(modrm2_not), .in2(modrm1_not), .in3(modrm0_not), .in4(op15_not), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not), .in11(op8), .in12(op7_not), .in13(op6_not), .in14(op5), .in15(op4_not), .in16(op3_not), .in17(op2_not), .in18(op1_not));
and16$ and_gate553(.out(and553), .in0(
sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8), .in9(op7_not), .in10(op6
), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and13$ and_gate554(.out(and554), .in0(modrm0_not), .in1(op15_not), .in2(op14), .in3(op13_not), .in4(op12), .in5(op11_not), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4));
and14$ and_gate555(.out(and555), .in0(sizeov_not), .in1(op13_not), .in2(op12), .in3(op11), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5_not), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate556(.out(and556), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op10_not), .in5(op9), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate557(.out(and557), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(op11_not), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7_not), .in8(op6), .in9(op5), .in10(op4_not), .in11(op3_not), .in12(op2), .in13(op1_not));
and14$ and_gate558(.out(and558), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4_not), .in5(op9_not), .in6(op8), .in7(op7), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and11$ and_gate559(.out(and559), .in0(modrm1_not), .in1(modrm0_not), .in2(op15_not), .in3(op14), .in4(op13_not), .in5(op12), .in6(op11_not), .in7(op10_not), .in8(op9), .in9(op8_not), .in10(op7));
and10$ and_gate560(.out(and560), .in0(modrm0), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op6_not), .in5(op5_not), .in6(op4_not), .in7(op3_not), .in8(op2_not), .in9(op1_not));
and8$ and_gate561(.out(and561), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(op11), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op1_not));
and8$ and_gate562(.out(and562), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7));
and8$ and_gate563(.out(and563), .in0(op14), .in1(op13), .in2(op12_not), .in3(op11_not), .in4(op4_not), .in5(op3_not), .in6(op2_not), .in7(op1_not));
and20$ and_gate564(.out(and564), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(modrm3), .in6(modrm2
), .in7(modrm1), .in8(modrm0), .in9(op15_not), .in10(op14_not), .in11(op13), .in12(op12_not), .in13(op11), .in14(op10), .in15(op9_not), .in16(op8_not), .in17(op7_not), .in18(op6
), .in19(op5));
and16$ and_gate565(.out(and565), .in0(sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5), .in4(modrm4_not), .in5(op11_not), .in6(op10_not), .in7(op9_not), .in8(op8
), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and13$ and_gate566(.out(and566), .in0(modrm0_not), .in1(op15_not), .in2(op14), .in3(op13_not), .in4(op12
), .in5(op11_not), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4));
and13$ and_gate567(.out(and567), .in0(sizeov_not), .in1(modrm7), .in2(modrm6
), .in3(modrm5), .in4(modrm4_not), .in5(modrm3_not), .in6(modrm2), .in7(modrm1_not), .in8(modrm0), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2));
and14$ and_gate568(.out(and568), .in0(
sizeov), .in1(modrm7_not), .in2(modrm6), .in3(modrm5_not), .in4(modrm4_not), .in5(modrm3_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate569(.out(and569), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(modrm4), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10), .in10(op9), .in11(op8), .in12(op7_not), .in13(op6));
and14$ and_gate570(.out(and570), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op10_not), .in5(op9), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5), .in10(op4), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate571(.out(and571), .in0(sizeov_not), .in1(modrm7_not), .in2(op12_not), .in3(op11), .in4(op10), .in5(op9_not), .in6(op8_not), .in7(op7), .in8(op6), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and14$ and_gate572(.out(and572), .in0(modrm4_not), .in1(modrm3_not), .in2(modrm2_not), .in3(modrm1_not), .in4(modrm0), .in5(op15), .in6(op14), .in7(op13_not), .in8(op12_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not));
and11$ and_gate573(.out(and573), .in0(modrm1_not), .in1(modrm0_not), .in2(op15_not), .in3(op14), .in4(op13_not), .in5(op12), .in6(op11_not), .in7(op10_not), .in8(op9), .in9(op8_not), .in10(op7));
and10$ and_gate574(.out(and574), .in0(sizeov), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5), .in4(modrm4_not), .in5(modrm3), .in6(op8
), .in7(op7), .in8(op6_not), .in9(op5));
and10$ and_gate575(.out(and575), .in0(modrm2_not), .in1(modrm1_not), .in2(modrm0_not), .in3(op15_not), .in4(op14_not), .in5(op13), .in6(op4_not), .in7(op3_not), .in8(op2), .in9(op1_not));
and9$ and_gate576(.out(and576), .in0(sizeov_not), .in1(modrm7_not), .in2(modrm6_not), .in3(modrm5_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9
), .in8(op8));
and8$ and_gate577(.out(and577), .in0(sizeov_not), .in1(modrm7), .in2(modrm6_not), .in3(modrm5), .in4(op10), .in5(op9), .in6(op8_not), .in7(op7));

or14$ or_gate0(.out(or0), .in0(and0), .in1(and1), .in2(and2), .in3(and3), .in4(and4), .in5(and5), .in6(and6), .in7(and7), .in8(and8), .in9(and9), .in10(and10), .in11(and11), .in12(and12), .in13(and13));
or12$ or_gate1(.out(or1), .in0(and14), .in1(and15), .in2(and16), .in3(and17), .in4(and18), .in5(and19), .in6(and20), .in7(and21), .in8(and22), .in9(and23), .in10(and24), .in11(and25));
or14$ or_gate2(.out(or2), .in0(and26), .in1(and27), .in2(and28), .in3(and29), .in4(and30), .in5(and31), .in6(and32), .in7(and33), .in8(and34), .in9(and35), .in10(and36), .in11(and37), .in12(and38), .in13(and39));
or8$ or_gate3(.out(or3), .in0(and40), .in1(and41), .in2(and42), .in3(and43), .in4(and44), .in5(and45), .in6(and46), .in7(and47));
or14$ or_gate4(.out(or4), .in0(and48), .in1(and49), .in2(and50), .in3(and51), .in4(and52), .in5(and53), .in6(and54), .in7(and55), .in8(and56), .in9(and57), .in10(and58), .in11(and59), .in12(and60), .in13(and61));
or18$ or_gate5(.out(or5), .in0(and62), .in1(and63), .in2(and64), .in3(and65), .in4(and66), .in5(and67), .in6(and68), .in7(and69), .in8(and70), .in9(and71), .in10(and72), .in11(and73), .in12(and74), .in13(and75), .in14(and76), .in15(and77), .in16(and78), .in17(and79));
or19$ or_gate6(.out(or6), .in0(and80), .in1(and81), .in2(and82), .in3(and83), .in4(and84), .in5(and85), .in6(and86), .in7(and87), .in8(and88), .in9(and89), .in10(and90), .in11(and91), .in12(and92), .in13(and93), .in14(and94), .in15(and95), .in16(and96), .in17(and97), .in18(and98));
or17$ or_gate7(.out(or7), .in0(and99), .in1(and100), .in2(and101), .in3(and102), .in4(and103), .in5(and104), .in6(and105), .in7(and106), .in8(and107), .in9(and108), .in10(and109), .in11(and110), .in12(and111), .in13(and112), .in14(and113), .in15(and114), .in16(and115));
or16$ or_gate8(.out(or8), .in0(and116), .in1(and117), .in2(and118), .in3(and119), .in4(and120), .in5(and121), .in6(and122), .in7(and123), .in8(and124), .in9(and125), .in10(and126), .in11(and127), .in12(and128), .in13(and129), .in14(and130), .in15(and131));
or14$ or_gate9(.out(or9), .in0(and132), .in1(and133), .in2(and134), .in3(and135), .in4(and136), .in5(and137), .in6(and138), .in7(and139), .in8(and140), .in9(and141), .in10(and142), .in11(and143), .in12(and144), .in13(and145));
or19$ or_gate10(.out(or10), .in0(and146), .in1(and147), .in2(and148), .in3(and149), .in4(and150), .in5(and151), .in6(and152), .in7(and153), .in8(and154), .in9(and155), .in10(and156), .in11(and157), .in12(and158), .in13(and159), .in14(and160), .in15(and161), .in16(and162), .in17(and163), .in18(and164));
or24$ or_gate11(.out(or11), .in0(and165), .in1(and166), .in2(and167), .in3(and168), .in4(and169), .in5(and170), .in6(and171), .in7(and172), .in8(and173), .in9(and174), .in10(and175), .in11(and176), .in12(and177), .in13(and178), .in14(and179), .in15(and180), .in16(and181), .in17(and182), .in18(and183), .in19(and184), .in20(and185), .in21(and186), .in22(and187), .in23(and188));
or26$ or_gate12(.out(or12), .in0(and189), .in1(and190), .in2(and191), .in3(and192), .in4(and193), .in5(and194), .in6(and195), .in7(and196), .in8(and197), .in9(and198), .in10(and199), .in11(and200), .in12(and201), .in13(and202), .in14(and203), .in15(and204), .in16(and205), .in17(and206), .in18(and207), .in19(and208), .in20(and209), .in21(and210), .in22(and211), .in23(and212), .in24(and213), .in25(and214));
or24$ or_gate13(.out(or13), .in0(and215), .in1(and216), .in2(and217), .in3(and218), .in4(and219), .in5(and220), .in6(and221), .in7(and222), .in8(and223), .in9(and224), .in10(and225), .in11(and226), .in12(and227), .in13(and228), .in14(and229), .in15(and230), .in16(and231), .in17(and232), .in18(and233), .in19(and234), .in20(and235), .in21(and236), .in22(and237), .in23(and238));
or23$ or_gate14(.out(or14), .in0(and239), .in1(and240), .in2(and241), .in3(and242), .in4(and243), .in5(and244), .in6(and245), .in7(and246), .in8(and247), .in9(and248), .in10(and249), .in11(and250), .in12(and251), .in13(and252), .in14(and253), .in15(and254), .in16(and255), .in17(and256), .in18(and257), .in19(and258), .in20(and259), .in21(and260), .in22(and261));
or20$ or_gate15(.out(or15), .in0(and262), .in1(and263), .in2(and264), .in3(and265), .in4(and266), .in5(and267), .in6(and268), .in7(and269), .in8(and270), .in9(and271), .in10(and272), .in11(and273), .in12(and274), .in13(and275), .in14(and276), .in15(and277), .in16(and278), .in17(and279), .in18(and280), .in19(and281));
or16$ or_gate16(.out(or16), .in0(and282), .in1(and283), .in2(and284), .in3(and285), .in4(and286), .in5(and287), .in6(and288), .in7(and289), .in8(and290), .in9(and291), .in10(and292), .in11(and293), .in12(and294), .in13(and295), .in14(and296), .in15(and297));
or22$ or_gate17(.out(or17), .in0(and298), .in1(and299), .in2(and300), .in3(and301), .in4(and302), .in5(and303), .in6(and304), .in7(and305), .in8(and306), .in9(and307), .in10(and308), .in11(and309), .in12(and310), .in13(and311), .in14(and312), .in15(and313), .in16(and314), .in17(and315), .in18(and316), .in19(and317), .in20(and318), .in21(and319));
or19$ or_gate18(.out(or18), .in0(and320), .in1(and321), .in2(and322), .in3(and323), .in4(and324), .in5(and325), .in6(and326), .in7(and327), .in8(and328), .in9(and329), .in10(and330), .in11(and331), .in12(and332), .in13(and333), .in14(and334), .in15(and335), .in16(and336), .in17(and337), .in18(and338));
or17$ or_gate19(.out(or19), .in0(and339), .in1(and340), .in2(and341), .in3(and342), .in4(and343), .in5(and344), .in6(and345), .in7(and346), .in8(and347), .in9(and348), .in10(and349), .in11(and350), .in12(and351), .in13(and352), .in14(and353), .in15(and354), .in16(and355));
or19$ or_gate20(.out(or20), .in0(and356), .in1(and357), .in2(and358), .in3(and359), .in4(and360), .in5(and361), .in6(and362), .in7(and363), .in8(and364), .in9(and365), .in10(and366), .in11(and367), .in12(and368), .in13(and369), .in14(and370), .in15(and371), .in16(and372), .in17(and373), .in18(and374));
or17$ or_gate21(.out(or21), .in0(and375), .in1(and376), .in2(and377), .in3(and378), .in4(and379), .in5(and380), .in6(and381), .in7(and382), .in8(and383), .in9(and384), .in10(and385), .in11(and386), .in12(and387), .in13(and388), .in14(and389), .in15(and390), .in16(and391));
or19$ or_gate22(.out(or22), .in0(and392), .in1(and393), .in2(and394), .in3(and395), .in4(and396), .in5(and397), .in6(and398), .in7(and399), .in8(and400), .in9(and401), .in10(and402), .in11(and403), .in12(and404), .in13(and405), .in14(and406), .in15(and407), .in16(and408), .in17(and409), .in18(and410));
or12$ or_gate23(.out(or23), .in0(and411), .in1(and412), .in2(and413), .in3(and414), .in4(and415), .in5(and416), .in6(and417), .in7(and418), .in8(and419), .in9(and420), .in10(and421), .in11(and422));
or12$ or_gate24(.out(or24), .in0(and423), .in1(and424), .in2(and425), .in3(and426), .in4(and427), .in5(and428), .in6(and429), .in7(and430), .in8(and431), .in9(and432), .in10(and433), .in11(and434));
or12$ or_gate25(.out(or25), .in0(and435), .in1(and436), .in2(and437), .in3(and438), .in4(and439), .in5(and440), .in6(and441), .in7(and442), .in8(and443), .in9(and444), .in10(and445), .in11(and446));
or10$ or_gate26(.out(or26), .in0(and447), .in1(and448), .in2(and449), .in3(and450), .in4(and451), .in5(and452), .in6(and453), .in7(and454), .in8(and455), .in9(and456));
or14$ or_gate27(.out(or27), .in0(and457), .in1(and458), .in2(and459), .in3(and460), .in4(and461), .in5(and462), .in6(and463), .in7(and464), .in8(and465), .in9(and466), .in10(and467), .in11(and468), .in12(and469), .in13(and470));
or18$ or_gate28(.out(or28), .in0(and471), .in1(and472), .in2(and473), .in3(and474), .in4(and475), .in5(and476), .in6(and477), .in7(and478), .in8(and479), .in9(and480), .in10(and481), .in11(and482), .in12(and483), .in13(and484), .in14(and485), .in15(and486), .in16(and487), .in17(and488));
or15$ or_gate29(.out(or29), .in0(and489), .in1(and490), .in2(and491), .in3(and492), .in4(and493), .in5(and494), .in6(and495), .in7(and496), .in8(and497), .in9(and498), .in10(and499), .in11(and500), .in12(and501), .in13(and502), .in14(and503));
or10$ or_gate30(.out(or30), .in0(and504), .in1(and505), .in2(and506), .in3(and507), .in4(and508), .in5(and509), .in6(and510), .in7(and511), .in8(and512), .in9(and513));
or11$ or_gate31(.out(or31), .in0(and514), .in1(and515), .in2(and516), .in3(and517), .in4(and518), .in5(and519), .in6(and520), .in7(and521), .in8(and522), .in9(and523), .in10(and524));
or11$ or_gate32(.out(or32), .in0(and525), .in1(and526), .in2(and527), .in3(and528), .in4(and529), .in5(and530), .in6(and531), .in7(and532), .in8(and533), .in9(and534), .in10(and535));
or13$ or_gate33(.out(or33), .in0(and536), .in1(and537), .in2(and538), .in3(and539), .in4(and540), .in5(and541), .in6(and542), .in7(and543), .in8(and544), .in9(and545), .in10(and546), .in11(and547), .in12(and548));
or15$ or_gate34(.out(or34), .in0(and549), .in1(and550), .in2(and551), .in3(and552), .in4(and553), .in5(and554), .in6(and555), .in7(and556), .in8(and557), .in9(and558), .in10(and559), .in11(and560), .in12(and561), .in13(and562), .in14(and563));
or14$ or_gate35(.out(or35), .in0(and564), .in1(and565), .in2(and566), .in3(and567), .in4(and568), .in5(and569), .in6(and570), .in7(and571), .in8(and572), .in9(and573), .in10(and574), .in11(and575), .in12(and576), .in13(and577));

assign setd = or0;
assign cleard = or1;
assign size2 = or2;
assign size1 = or3;
assign size0 = or4;
assign op0_2 = or5;
assign op0_1 = or6;
assign op0_0 = or7;
assign op1_2 = or8;
assign op1_1 = or9;
assign op1_0 = or10;
assign op0_reg_4 = or11;
assign op0_reg_3 = or12;
assign op0_reg_2 = or13;
assign op0_reg_1 = or14;
assign op0_reg_0 = or15;
assign op1_reg_4 = or16;
assign op1_reg_3 = or17;
assign op1_reg_2 = or18;
assign op1_reg_1 = or19;
assign op1_reg_0 = or20;
assign alu_op_3 = or21;
assign alu_op_2 = or22;
assign alu_op_1 = or23;
assign alu_op_0 = or24;
assign flag0_2 = or25;
assign flag0_1 = or26;
assign flag0_0 = or27;
assign flag1_2 = or28;
assign flag1_1 = or29;
assign flag1_0 = or30;
assign stack_op_1 = or31;
assign stack_op_0 = or32;
assign rom_control_2 = or33;
assign rom_control_1 = or34;
assign rom_control_0 = or35;
endmodule
