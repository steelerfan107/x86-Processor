module dcache();

endmodule
