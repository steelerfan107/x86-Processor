module mem_align(
    input [31:0] reg_out,
    input [1:0] wr_size,
    input [31:0] mem_data,
    input [1:0] off,
    output [31:0] out
);

    

endmodule
