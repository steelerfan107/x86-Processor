module opcode_modrm_control_cloud (
 input  sizeov,				    
 input 	modrm7, 
 input 	modrm6, 
 input 	modrm5, 
 input 	modrm4, 
 input 	modrm3, 
 input 	modrm2, 
 input 	modrm1, 
 input 	modrm0, 
 input 	op15, 
 input 	op14, 
 input 	op13, 
 input 	op12, 
 input 	op11, 
 input 	op10, 
 input 	op9, 
 input 	op8, 
 input 	op7, 
 input 	op6, 
 input 	op5, 
 input 	op4, 
 input 	op3, 
 input 	op2, 
 input 	op1, 
 input 	op0,
 output setd, 
 output cleard, 
 output size2, 
 output size1, 
 output size0, 
 output op0_2, 
 output op0_1, 
 output op0_0, 
 output op1_2, 
 output op1_1, 
 output op1_0, 
 output op0_reg_4, 
 output op0_reg_3, 
 output op0_reg_2, 
 output op0_reg_1, 
 output op0_reg_0, 
 output op1_reg_4, 
 output op1_reg_3, 
 output op1_reg_2, 
 output op1_reg_1, 
 output op1_reg_0, 
 output alu_op_3, 
 output alu_op_2, 
 output alu_op_1, 
 output alu_op_0, 
 output flag0_2, 
 output flag0_1, 
 output flag0_0, 
 output flag1_2, 
 output flag1_1, 
 output flag1_0, 
 output stack_op_1, 
 output stack_op_0				   
);

wire sizeov_not;
wire op9_not;
wire op7_not;
wire op6_not;
wire op5_not;
wire op4_not;
wire op3_not;
wire op2_not;
wire op1_not;
wire op0_not;
wire and0;
wire op8_not;
wire op5_not;
wire op4_not;
wire and1;
wire op15_not;
wire op14_not;
wire op13_not;
wire op12_not;
wire and2;
wire and3;
wire op14_not;
wire and4;
wire sizeov_not;
wire and5;
wire and6;
wire op10_not;
wire and7;
wire or0;
wire and8;
wire op10_not;
wire op6_not;
wire and9;
wire and10;
wire op15_not;
wire and11;
wire and12;
wire op11_not;
wire and13;
wire op12_not;
wire and14;
wire sizeov_not;
wire op2_not;
wire and15;
wire op7_not;
wire and16;
wire and17;
wire op15_not;
wire op3_not;
wire and18;
wire and19;
wire op13_not;
wire and20;
wire and21;
wire and22;
wire and23;
wire and24;
wire and25;
wire and26;
wire modrm5_not;
wire modrm3_not;
wire and27;
wire op11_not;
wire and28;
wire and29;
wire and30;
wire modrm3_not;
wire and31;
wire op9_not;
wire and32;
wire modrm4_not;
wire and33;
wire op1_not;
wire and34;
wire and35;
wire and36;
wire and37;
wire modrm5_not;
wire and38;
wire and39;
wire and40;
wire and41;
wire and42;
wire and43;
wire and44;
wire modrm5_not;
wire and45;
wire and46;
wire and47;
wire and48;
wire and49;
wire and50;
wire or1;
wire and51;
wire and52;
wire and53;
wire and54;
wire and55;
wire and56;
wire and57;
wire and58;
wire and59;
wire and60;
wire and61;
wire and62;
wire and63;
wire and64;
wire and65;
wire and66;
wire and67;
wire and68;
wire and69;
wire and70;
wire and71;
wire and72;
wire and73;
wire and74;
wire and75;
wire and76;
wire and77;
wire and78;
wire and79;
wire and80;
wire and81;
wire modrm4_not;
wire and82;
wire and83;
wire and84;
wire and85;
wire and86;
wire and87;
wire or2;
wire and88;
wire op8_not;
wire and89;
wire and90;
wire and91;
wire and92;
wire and93;
wire and94;
wire and95;
wire and96;
wire and97;
wire and98;
wire and99;
wire and100;
wire and101;
wire and102;
wire and103;
wire and104;
wire and105;
wire and106;
wire and107;
wire and108;
wire and109;
wire and110;
wire and111;
wire and112;
wire and113;
wire and114;
wire and115;
wire and116;
wire and117;
wire and118;
wire and119;
wire and120;
wire and121;
wire and122;
wire and123;
wire and124;
wire or3;
wire and125;
wire and126;
wire and127;
wire and128;
wire and129;
wire and130;
wire and131;
wire and132;
wire and133;
wire or4;
wire and134;
wire and135;
wire and136;
wire and137;
wire and138;
wire and139;
wire and140;
wire and141;
wire and142;
wire and143;
wire and144;
wire and145;
wire and146;
wire and147;
wire and148;
wire and149;
wire and150;
wire and151;
wire and152;
wire and153;
wire and154;
wire and155;
wire and156;
wire and157;
wire and158;
wire and159;
wire or5;
wire and160;
wire and161;
wire and162;
wire and163;
wire and164;
wire and165;
wire and166;
wire and167;
wire and168;
wire and169;
wire and170;
wire and171;
wire and172;
wire and173;
wire and174;
wire and175;
wire and176;
wire and177;
wire and178;
wire and179;
wire and180;
wire and181;
wire and182;
wire and183;
wire and184;
wire and185;
wire and186;
wire and187;
wire and188;
wire and189;
wire and190;
wire and191;
wire and192;
wire and193;
wire and194;
wire and195;
wire or6;
wire and196;
wire and197;
wire and198;
wire and199;
wire and200;
wire and201;
wire or7;
wire and202;
wire and203;
wire and204;
wire and205;
wire and206;
wire and207;
wire and208;
wire and209;
wire and210;
wire and211;
wire and212;
wire and213;
wire and214;
wire and215;
wire and216;
wire and217;
wire and218;
wire and219;
wire and220;
wire and221;
wire and222;
wire and223;
wire and224;
wire and225;
wire and226;
wire and227;
wire and228;
wire and229;
wire and230;
wire and231;
wire and232;
wire and233;
wire and234;
wire and235;
wire and236;
wire or8;
wire and237;
wire and238;
wire or9;
wire and239;
wire and240;
wire and241;
wire and242;
wire and243;
wire and244;
wire and245;
wire and246;
wire and247;
wire and248;
wire and249;
wire and250;
wire and251;
wire and252;
wire and253;
wire or10;
wire and254;
wire and255;
wire or11;
wire and256;
wire and257;
wire and258;
wire or12;
wire and259;
wire and260;
wire and261;
wire or13;
wire and262;
wire and263;
wire and264;
wire and265;
wire and266;
wire and267;
wire and268;
wire and269;
wire and270;
wire and271;
wire and272;
wire or14;
wire and273;
wire and274;
wire and275;
wire and276;
wire or15;
wire and277;
wire and278;
wire and279;
wire and280;
wire and281;
wire and282;
wire and283;
wire and284;
wire and285;
wire and286;
wire and287;
wire and288;
wire and289;
wire and290;
wire and291;
wire and292;
wire and293;
wire and294;
wire and295;
wire and296;
wire or16;
wire and297;
wire and298;
wire and299;
wire and300;
wire and301;
wire and302;
wire and303;
wire and304;
wire and305;
wire and306;
wire and307;
wire and308;
wire and309;
wire and310;
wire and311;
wire and312;
wire and313;
wire and314;
wire and315;
wire and316;
wire and317;
wire and318;
wire and319;
wire and320;
wire and321;
wire and322;
wire and323;
wire and324;
wire and325;
wire and326;
wire and327;
wire and328;
wire and329;
wire and330;
wire and331;
wire and332;
wire and333;
wire and334;
wire and335;
wire and336;
wire and337;
wire and338;
wire and339;
wire and340;
wire or17;
wire and341;
wire and342;
wire and343;
wire and344;
wire and345;
wire and346;
wire and347;
wire and348;
wire and349;
wire and350;
wire and351;
wire and352;
wire and353;
wire and354;
wire and355;
wire and356;
wire and357;
wire and358;
wire and359;
wire and360;
wire and361;
wire or18;
wire and362;
wire and363;
wire and364;
wire and365;
wire and366;
wire and367;
wire and368;
wire and369;
wire and370;
wire and371;
wire and372;
wire and373;
wire and374;
wire and375;
wire and376;
wire and377;
wire or19;
wire and378;
wire and379;
wire and380;
wire and381;
wire or20;
wire and382;
wire and383;
wire and384;
wire or21;
wire and385;
wire and386;
wire or22;
wire and387;
wire and388;
wire and389;
wire and390;
wire and391;
wire and392;
wire or23;
wire and393;
wire and394;
wire and395;
wire and396;
wire and397;
wire and398;
wire and399;
wire or24;

inv1$ sizeov_inv (.out(sizeov_not), .in(sizeov));
inv1$ op9_inv (.out(op9_not), .in(op9));
inv1$ op7_inv (.out(op7_not), .in(op7));
inv1$ op6_inv (.out(op6_not), .in(op6));
inv1$ op5_inv (.out(op5_not), .in(op5));
inv1$ op4_inv (.out(op4_not), .in(op4));
inv1$ op3_inv (.out(op3_not), .in(op3));
inv1$ op2_inv (.out(op2_not), .in(op2));
inv1$ op1_inv (.out(op1_not), .in(op1));
inv1$ op0_inv (.out(op0_not), .in(op0));
inv1$ op8_inv (.out(op8_not), .in(op8));
inv1$ op15_inv (.out(op15_not), .in(op15));
inv1$ op14_inv (.out(op14_not), .in(op14));
inv1$ op13_inv (.out(op13_not), .in(op13));
inv1$ op12_inv (.out(op12_not), .in(op12));
inv1$ op10_inv (.out(op10_not), .in(op10));
inv1$ op11_inv (.out(op11_not), .in(op11));
inv1$ modrm5_inv (.out(modrm5_not), .in(modrm5));
inv1$ modrm3_inv (.out(modrm3_not), .in(modrm3));
inv1$ modrm4_inv (.out(modrm4_not), .in(modrm4));

and17$ and_gate0(.out(and0), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13), .in4(op12), .in5(op11), .in6(op10), .in7(op9_not), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and17$ and_gate1(.out(and1), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13), .in4(op12), .in5(op11), .in6(op10), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and17$ and_gate2(.out(and2), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5
), .in12(op4), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and17$ and_gate3(.out(and3), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10
), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not), .in16(op0));
and17$ and_gate4(.out(and4), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and16$ and_gate5(.out(and5), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op3), .in13(op2
), .in14(op1), .in15(op0_not));
and16$ and_gate6(.out(and6), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7
), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op1), .in15(op0_not));
and17$ and_gate7(.out(and7), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate8(.out(and8), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3
), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate9(.out(and9), .in0(op15), .in1(op14), .in2(op13), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate10(.out(and10), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13_not), .in4(op12_not), .in5(op10_not), .in6(op9), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate11(.out(and11), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and17$ and_gate12(.out(and12), .in0(
sizeov), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate13(.out(and13), .in0(sizeov_not), .in1(op14_not), .in2(op13), .in3(op12_not), .in4(op11_not), .in5(op10), .in6(op9_not), .in7(op8
), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate14(.out(and14), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and17$ and_gate15(.out(and15), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and17$ and_gate16(.out(and16), .in0(sizeov), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and17$ and_gate17(.out(and17), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate18(.out(and18), .in0(op15_not), .in1(op14), .in2(op13), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate19(.out(and19), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10), .in7(op9), .in8(op8
), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate20(.out(and20), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate21(.out(and21), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate22(.out(and22), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op11_not), .in5(op10), .in6(op9), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate23(.out(and23), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1), .in16(op0_not));
and15$ and_gate24(.out(and24), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate25(.out(and25), .in0(op15_not), .in1(op14_not), .in2(op13), .in3(op12_not), .in4(op11_not), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate26(.out(and26), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op9_not), .in6(op8
), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and10$ and_gate27(.out(and27), .in0(modrm5_not), .in1(modrm4), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13), .in6(op12), .in7(op10), .in8(op9), .in9(op8));
and16$ and_gate28(.out(and28), .in0(op15_not), .in1(op14_not), .in2(op13), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate29(.out(and29), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2), .in15(op0));
and16$ and_gate30(.out(and30), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op11_not), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate31(.out(and31), .in0(modrm5), .in1(modrm4), .in2(modrm3_not), .in3(op15), .in4(op14
), .in5(op13), .in6(op12), .in7(op11), .in8(op10), .in9(op9), .in10(op8));
and15$ and_gate32(.out(and32), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and12$ and_gate33(.out(and33), .in0(sizeov_not), .in1(modrm5
), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13), .in7(op12), .in8(op11), .in9(op10), .in10(op9), .in11(op8));
and16$ and_gate34(.out(and34), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate35(.out(and35), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and15$ and_gate36(.out(and36), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op8
), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate37(.out(and37), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate38(.out(and38), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11), .in8(op10), .in9(op9), .in10(op8));
and10$ and_gate39(.out(and39), .in0(
modrm5), .in1(modrm4), .in2(modrm3), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate40(.out(and40), .in0(modrm5
), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11_not), .in8(op10_not), .in9(op8));
and11$ and_gate41(.out(and41), .in0(modrm5
), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not), .in10(op8));
and11$ and_gate42(.out(and42), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op9), .in10(op8));
and10$ and_gate43(.out(and43), .in0(
modrm5), .in1(modrm4), .in2(modrm3), .in3(op15), .in4(op14), .in5(op13_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate44(.out(and44), .in0(modrm5
), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate45(.out(and45), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate46(.out(and46), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op8));
and11$ and_gate47(.out(and47), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op8));
and5$ and_gate48(.out(and48), .in0(op15_not), .in1(op14), .in2(op13_not), .in3(op12), .in4(op11));
and5$ and_gate49(.out(and49), .in0(op15), .in1(op14_not), .in2(op13), .in3(op12), .in4(op11));
and5$ and_gate50(.out(and50), .in0(op15
), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and17$ and_gate51(.out(and51), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5
), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not), .in16(op0_not));
and17$ and_gate52(.out(and52), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10
), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5), .in12(op4), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and17$ and_gate53(.out(and53), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not), .in16(op0));
and17$ and_gate54(.out(and54), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and16$ and_gate55(.out(and55), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9
), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op3), .in13(op2), .in14(op1), .in15(op0_not));
and16$ and_gate56(.out(and56), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op1), .in15(op0_not));
and15$ and_gate57(.out(and57), .in0(sizeov_not), .in1(op14
), .in2(op13), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op8_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and17$ and_gate58(.out(and58), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate59(.out(and59), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10
), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate60(.out(and60), .in0(sizeov_not), .in1(op15_not), .in2(op14), .in3(op13
), .in4(op12), .in5(op11_not), .in6(op10), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate61(.out(and61), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate62(.out(and62), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8
), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1), .in16(op0_not));
and15$ and_gate63(.out(and63), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13
), .in4(op12_not), .in5(op11_not), .in6(op9_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate64(.out(and64), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate65(.out(and65), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7
), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2), .in15(op0));
and10$ and_gate66(.out(and66), .in0(sizeov_not), .in1(modrm4), .in2(modrm3_not), .in3(op15), .in4(op13
), .in5(op12), .in6(op11), .in7(op10), .in8(op9), .in9(op8));
and11$ and_gate67(.out(and67), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4), .in3(modrm3_not), .in4(op15), .in5(op14
), .in6(op13), .in7(op12), .in8(op11_not), .in9(op10), .in10(op9));
and12$ and_gate68(.out(and68), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15
), .in5(op14), .in6(op13), .in7(op12), .in8(op11), .in9(op10), .in10(op9), .in11(op8));
and11$ and_gate69(.out(and69), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op11), .in8(op10), .in9(op9), .in10(op8));
and15$ and_gate70(.out(and70), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op9_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate71(.out(and71), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and14$ and_gate72(.out(and72), .in0(sizeov_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op7_not), .in7(op6_not), .in8(op5_not), .in9(op4_not), .in10(op3_not), .in11(op2_not), .in12(op1_not), .in13(op0_not));
and16$ and_gate73(.out(and73), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate74(.out(and74), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and10$ and_gate75(.out(and75), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op8));
and16$ and_gate76(.out(and76), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate77(.out(and77), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and11$ and_gate78(.out(and78), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and10$ and_gate79(.out(and79), .in0(sizeov_not), .in1(modrm5), .in2(modrm4), .in3(modrm3), .in4(op15
), .in5(op14), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op10_not));
and10$ and_gate80(.out(and80), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15
), .in5(op14), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op10_not));
and11$ and_gate81(.out(and81), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15
), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and11$ and_gate82(.out(and82), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10), .in10(op9));
and10$ and_gate83(.out(and83), .in0(sizeov_not), .in1(modrm5
), .in2(modrm4), .in3(modrm3), .in4(op15), .in5(op14), .in6(op13_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate84(.out(and84), .in0(sizeov_not), .in1(modrm5
), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and11$ and_gate85(.out(and85), .in0(sizeov_not), .in1(modrm5
), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op8));
and6$ and_gate86(.out(and86), .in0(sizeov_not), .in1(op15_not), .in2(op14), .in3(op13_not), .in4(op12), .in5(op11));
and5$ and_gate87(.out(and87), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op12), .in4(op11));
and17$ and_gate88(.out(and88), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5
), .in12(op4), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and16$ and_gate89(.out(and89), .in0(op15), .in1(op14), .in2(op13), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate90(.out(and90), .in0(sizeov), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate91(.out(and91), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and17$ and_gate92(.out(and92), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate93(.out(and93), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and15$ and_gate94(.out(and94), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate95(.out(and95), .in0(sizeov_not), .in1(op15_not), .in2(op14), .in3(op13), .in4(op12), .in5(op11_not), .in6(op10), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate96(.out(and96), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate97(.out(and97), .in0(sizeov_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and15$ and_gate98(.out(and98), .in0(op15_not), .in1(op14_not), .in2(op12_not), .in3(op11_not), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and10$ and_gate99(.out(and99), .in0(modrm5_not), .in1(modrm4), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13), .in6(op12
), .in7(op10), .in8(op9), .in9(op8));
and16$ and_gate100(.out(and100), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8
), .in9(op7), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2), .in15(op0));
and15$ and_gate101(.out(and101), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and11$ and_gate102(.out(and102), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13), .in7(op12), .in8(op11_not), .in9(op10), .in10(op9));
and12$ and_gate103(.out(and103), .in0(sizeov_not), .in1(modrm5
), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13), .in7(op12), .in8(op11), .in9(op10), .in10(op9), .in11(op8));
and16$ and_gate104(.out(and104), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate105(.out(and105), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate106(.out(and106), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate107(.out(and107), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and11$ and_gate108(.out(and108), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11), .in8(op10), .in9(op9), .in10(op8));
and11$ and_gate109(.out(and109), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and10$ and_gate110(.out(and110), .in0(modrm5), .in1(modrm4), .in2(modrm3), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate111(.out(and111), .in0(sizeov_not), .in1(modrm5), .in2(modrm4), .in3(modrm3), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op10_not));
and10$ and_gate112(.out(and112), .in0(
modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate113(.out(and113), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op10_not));
and11$ and_gate114(.out(and114), .in0(
modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not), .in10(op8));
and11$ and_gate115(.out(and115), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and11$ and_gate116(.out(and116), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op9), .in10(op8));
and11$ and_gate117(.out(and117), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10), .in10(op9));
and10$ and_gate118(.out(and118), .in0(
modrm5), .in1(modrm4), .in2(modrm3), .in3(op15), .in4(op14), .in5(op13_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate119(.out(and119), .in0(sizeov_not), .in1(modrm5), .in2(modrm4), .in3(modrm3), .in4(op15), .in5(op14), .in6(op13_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate120(.out(and120), .in0(modrm5
), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate121(.out(and121), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate122(.out(and122), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate123(.out(and123), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op8));
and11$ and_gate124(.out(and124), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op8));
and17$ and_gate125(.out(and125), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5
), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not), .in16(op0));
and17$ and_gate126(.out(and126), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10
), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and16$ and_gate127(.out(and127), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op3), .in13(op2), .in14(op1), .in15(op0_not));
and16$ and_gate128(.out(and128), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op1), .in15(op0_not));
and16$ and_gate129(.out(and129), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8
), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and17$ and_gate130(.out(and130), .in0(sizeov), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and17$ and_gate131(.out(and131), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate132(.out(and132), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate133(.out(and133), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op11_not), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate134(.out(and134), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5
), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not), .in16(op0));
and17$ and_gate135(.out(and135), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10
), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and16$ and_gate136(.out(and136), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op3), .in13(op2), .in14(op1), .in15(op0_not));
and16$ and_gate137(.out(and137), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate138(.out(and138), .in0(op15), .in1(op14), .in2(op13), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate139(.out(and139), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11
), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op1), .in15(op0_not));
and17$ and_gate140(.out(and140), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and17$ and_gate141(.out(and141), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate142(.out(and142), .in0(sizeov_not), .in1(op15_not), .in2(op14), .in3(op13), .in4(op12), .in5(op11_not), .in6(op10), .in7(op8
), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate143(.out(and143), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and15$ and_gate144(.out(and144), .in0(op15_not), .in1(op14_not), .in2(op12_not), .in3(op11_not), .in4(op10), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and17$ and_gate145(.out(and145), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1), .in16(op0_not));
and15$ and_gate146(.out(and146), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op12_not), .in4(op11_not), .in5(op10), .in6(op9_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate147(.out(and147), .in0(op15_not), .in1(op14_not), .in2(op13), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate148(.out(and148), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate149(.out(and149), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2), .in15(op0));
and15$ and_gate150(.out(and150), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11), .in4(op10_not), .in5(op9), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate151(.out(and151), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate152(.out(and152), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate153(.out(and153), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and15$ and_gate154(.out(and154), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op10), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate155(.out(and155), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate156(.out(and156), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and5$ and_gate157(.out(and157), .in0(op15_not), .in1(op14), .in2(op13_not), .in3(op12), .in4(op11));
and5$ and_gate158(.out(and158), .in0(op15), .in1(op14_not), .in2(op13), .in3(op12), .in4(op11));
and5$ and_gate159(.out(and159), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and17$ and_gate160(.out(and160), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5
), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not), .in16(op0));
and17$ and_gate161(.out(and161), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10
), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and16$ and_gate162(.out(and162), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op3), .in13(op2), .in14(op1), .in15(op0_not));
and16$ and_gate163(.out(and163), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate164(.out(and164), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6
), .in11(op5), .in12(op4_not), .in13(op3), .in14(op1), .in15(op0_not));
and16$ and_gate165(.out(and165), .in0(sizeov_not), .in1(op15_not), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate166(.out(and166), .in0(sizeov), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate167(.out(and167), .in0(op15_not), .in1(op14), .in2(op13), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate168(.out(and168), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11
), .in6(op10_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate169(.out(and169), .in0(sizeov_not), .in1(op15
), .in2(op14_not), .in3(op13), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and15$ and_gate170(.out(and170), .in0(op15_not), .in1(op14_not), .in2(op12_not), .in3(op11_not), .in4(op10), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and17$ and_gate171(.out(and171), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10
), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1), .in16(op0_not));
and15$ and_gate172(.out(and172), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op12_not), .in4(op11_not), .in5(op10), .in6(op9_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate173(.out(and173), .in0(op15_not), .in1(op14_not), .in2(op13), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate174(.out(and174), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9
), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate175(.out(and175), .in0(modrm5), .in1(modrm4), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13), .in6(op12), .in7(op11), .in8(op10), .in9(op9), .in10(op8));
and15$ and_gate176(.out(and176), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11
), .in4(op10_not), .in5(op9), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate177(.out(and177), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate178(.out(and178), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate179(.out(and179), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and15$ and_gate180(.out(and180), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op10), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate181(.out(and181), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate182(.out(and182), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3
), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and11$ and_gate183(.out(and183), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and11$ and_gate184(.out(and184), .in0(modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not), .in10(op8));
and11$ and_gate185(.out(and185), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and11$ and_gate186(.out(and186), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op9), .in10(op8));
and11$ and_gate187(.out(and187), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10), .in10(op9));
and10$ and_gate188(.out(and188), .in0(
modrm5), .in1(modrm4), .in2(modrm3), .in3(op15), .in4(op14), .in5(op13_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate189(.out(and189), .in0(sizeov_not), .in1(modrm5), .in2(modrm4), .in3(modrm3), .in4(op15), .in5(op14), .in6(op13_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate190(.out(and190), .in0(modrm5
), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate191(.out(and191), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate192(.out(and192), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate193(.out(and193), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op8));
and11$ and_gate194(.out(and194), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op8));
and5$ and_gate195(.out(and195), .in0(
op15), .in1(op14_not), .in2(op13), .in3(op12), .in4(op11));
and17$ and_gate196(.out(and196), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5
), .in12(op4), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and17$ and_gate197(.out(and197), .in0(sizeov), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate198(.out(and198), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate199(.out(and199), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate200(.out(and200), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op11_not), .in5(op10), .in6(op9), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate201(.out(and201), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13
), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate202(.out(and202), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5
), .in12(op4), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and16$ and_gate203(.out(and203), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8
), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and16$ and_gate204(.out(and204), .in0(sizeov_not), .in1(op15_not), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate205(.out(and205), .in0(op15_not), .in1(op14), .in2(op13), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate206(.out(and206), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7
), .in10(op6_not), .in11(op5), .in12(op4), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate207(.out(and207), .in0(sizeov_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and15$ and_gate208(.out(and208), .in0(op15_not), .in1(op14_not), .in2(op12_not), .in3(op11_not), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate209(.out(and209), .in0(op15_not), .in1(op14_not), .in2(op13), .in3(op12_not), .in4(op11_not), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate210(.out(and210), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13), .in4(op12_not), .in5(op11_not), .in6(op9_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate211(.out(and211), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate212(.out(and212), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op9_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate213(.out(and213), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op10), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate214(.out(and214), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate215(.out(and215), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate216(.out(and216), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate217(.out(and217), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and11$ and_gate218(.out(and218), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and10$ and_gate219(.out(and219), .in0(modrm5), .in1(modrm4), .in2(modrm3), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12
), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate220(.out(and220), .in0(sizeov_not), .in1(modrm5), .in2(modrm4), .in3(modrm3), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op10_not));
and10$ and_gate221(.out(and221), .in0(modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12
), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate222(.out(and222), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op10_not));
and11$ and_gate223(.out(and223), .in0(modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not), .in10(op8));
and11$ and_gate224(.out(and224), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and11$ and_gate225(.out(and225), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14
), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op9), .in10(op8));
and11$ and_gate226(.out(and226), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10), .in10(op9));
and10$ and_gate227(.out(and227), .in0(modrm5), .in1(modrm4), .in2(modrm3), .in3(op15
), .in4(op14), .in5(op13_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate228(.out(and228), .in0(sizeov_not), .in1(modrm5), .in2(modrm4), .in3(modrm3
), .in4(op15), .in5(op14), .in6(op13_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate229(.out(and229), .in0(modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(op15
), .in4(op14), .in5(op13_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate230(.out(and230), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate231(.out(and231), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3), .in3(op15
), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate232(.out(and232), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15
), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op8));
and11$ and_gate233(.out(and233), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op8));
and5$ and_gate234(.out(and234), .in0(op15_not), .in1(op14), .in2(op13_not), .in3(op12
), .in4(op11));
and5$ and_gate235(.out(and235), .in0(op15), .in1(op14_not), .in2(op13), .in3(op12), .in4(op11));
and5$ and_gate236(.out(and236), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and5$ and_gate237(.out(and237), .in0(op15_not), .in1(op14), .in2(op13_not), .in3(op12), .in4(op11));
and5$ and_gate238(.out(and238), .in0(op15), .in1(op14_not), .in2(op13), .in3(op12), .in4(op11));
and17$ and_gate239(.out(and239), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6
), .in11(op5), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not), .in16(op0));
and17$ and_gate240(.out(and240), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11
), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and16$ and_gate241(.out(and241), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op3), .in13(op2), .in14(op1), .in15(op0_not));
and16$ and_gate242(.out(and242), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3), .in13(op2
), .in14(op1_not), .in15(op0_not));
and16$ and_gate243(.out(and243), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7
), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op1), .in15(op0_not));
and17$ and_gate244(.out(and244), .in0(sizeov), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11
), .in6(op10), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate245(.out(and245), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate246(.out(and246), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1), .in16(op0_not));
and15$ and_gate247(.out(and247), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11
), .in5(op10_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate248(.out(and248), .in0(op15_not), .in1(op14_not), .in2(op13), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate249(.out(and249), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate250(.out(and250), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate251(.out(and251), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate252(.out(and252), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and15$ and_gate253(.out(and253), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11
), .in5(op10_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate254(.out(and254), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and16$ and_gate255(.out(and255), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10
), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate256(.out(and256), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11_not), .in6(op10), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate257(.out(and257), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11
), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and17$ and_gate258(.out(and258), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate259(.out(and259), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2_not), .in15(op1_not));
and17$ and_gate260(.out(and260), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10
), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and17$ and_gate261(.out(and261), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and5$ and_gate262(.out(and262), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and17$ and_gate263(.out(and263), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6
), .in11(op5), .in12(op4), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and17$ and_gate264(.out(and264), .in0(sizeov), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10
), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate265(.out(and265), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and16$ and_gate266(.out(and266), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4
), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and15$ and_gate267(.out(and267), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate268(.out(and268), .in0(sizeov_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and15$ and_gate269(.out(and269), .in0(op15_not), .in1(op14_not), .in2(op12_not), .in3(op11_not), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate270(.out(and270), .in0(op14_not), .in1(op13_not), .in2(op12_not), .in3(op11), .in4(op10_not), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate271(.out(and271), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10), .in6(op9
), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate272(.out(and272), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and10$ and_gate273(.out(and273), .in0(modrm5), .in1(modrm4), .in2(modrm3), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate274(.out(and274), .in0(sizeov_not), .in1(modrm5), .in2(modrm4), .in3(modrm3), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op10_not));
and10$ and_gate275(.out(and275), .in0(
modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate276(.out(and276), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op10_not));
and17$ and_gate277(.out(and277), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5
), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not), .in16(op0));
and16$ and_gate278(.out(and278), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10
), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op3), .in13(op2), .in14(op1), .in15(op0_not));
and16$ and_gate279(.out(and279), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op1), .in15(op0_not));
and16$ and_gate280(.out(and280), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and15$ and_gate281(.out(and281), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate282(.out(and282), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op9_not), .in6(op8
), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate283(.out(and283), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate284(.out(and284), .in0(
op15), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate285(.out(and285), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate286(.out(and286), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and10$ and_gate287(.out(and287), .in0(modrm5), .in1(modrm4
), .in2(modrm3), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate288(.out(and288), .in0(sizeov_not), .in1(modrm5
), .in2(modrm4), .in3(modrm3), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op10_not));
and10$ and_gate289(.out(and289), .in0(modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate290(.out(and290), .in0(sizeov_not), .in1(modrm5
), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op10_not));
and10$ and_gate291(.out(and291), .in0(modrm5), .in1(modrm4
), .in2(modrm3), .in3(op15), .in4(op14), .in5(op13_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate292(.out(and292), .in0(sizeov_not), .in1(modrm5
), .in2(modrm4), .in3(modrm3), .in4(op15), .in5(op14), .in6(op13_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate293(.out(and293), .in0(modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate294(.out(and294), .in0(sizeov_not), .in1(modrm5
), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate295(.out(and295), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op8));
and5$ and_gate296(.out(and296), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and17$ and_gate297(.out(and297), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6
), .in11(op5), .in12(op4), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and17$ and_gate298(.out(and298), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11
), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op2), .in15(op1), .in16(op0));
and16$ and_gate299(.out(and299), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and17$ and_gate300(.out(and300), .in0(
sizeov), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9_not), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate301(.out(and301), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8
), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and17$ and_gate302(.out(and302), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13
), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate303(.out(and303), .in0(sizeov_not), .in1(op15_not), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate304(.out(and304), .in0(sizeov), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and17$ and_gate305(.out(and305), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13
), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate306(.out(and306), .in0(op15_not), .in1(op14), .in2(op13), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate307(.out(and307), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10), .in7(op9), .in8(op8
), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate308(.out(and308), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate309(.out(and309), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and11$ and_gate310(.out(and310), .in0(modrm5_not), .in1(modrm4), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13), .in6(op12), .in7(op11_not), .in8(op10), .in9(op9), .in10(op8));
and16$ and_gate311(.out(and311), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8
), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate312(.out(and312), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op11_not), .in5(op10), .in6(op9), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate313(.out(and313), .in0(sizeov_not), .in1(op15_not), .in2(op14), .in3(op13), .in4(op12), .in5(op11_not), .in6(op10), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate314(.out(and314), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1), .in16(op0_not));
and16$ and_gate315(.out(and315), .in0(sizeov_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11
), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and15$ and_gate316(.out(and316), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13_not), .in4(op12_not), .in5(op10_not), .in6(op9), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate317(.out(and317), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2), .in15(op0));
and16$ and_gate318(.out(and318), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op11_not), .in5(op10), .in6(op9
), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate319(.out(and319), .in0(modrm5), .in1(modrm4), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13), .in6(op12), .in7(op11), .in8(op10), .in9(op9), .in10(op8));
and11$ and_gate320(.out(and320), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4
), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13), .in7(op12), .in8(op11_not), .in9(op10), .in10(op9));
and12$ and_gate321(.out(and321), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13), .in7(op12), .in8(op11), .in9(op10), .in10(op9), .in11(op8));
and16$ and_gate322(.out(and322), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate323(.out(and323), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and15$ and_gate324(.out(and324), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate325(.out(and325), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10
), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate326(.out(and326), .in0(sizeov_not), .in1(op15
), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate327(.out(and327), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11), .in8(op10
), .in9(op9), .in10(op8));
and10$ and_gate328(.out(and328), .in0(modrm5), .in1(modrm4), .in2(modrm3), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate329(.out(and329), .in0(sizeov_not), .in1(modrm5), .in2(modrm4), .in3(modrm3), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op10_not));
and10$ and_gate330(.out(and330), .in0(
modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate331(.out(and331), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op10_not));
and11$ and_gate332(.out(and332), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10), .in9(op9), .in10(op8));
and11$ and_gate333(.out(and333), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10), .in10(op9));
and10$ and_gate334(.out(and334), .in0(
modrm5), .in1(modrm4), .in2(modrm3), .in3(op15), .in4(op14), .in5(op13_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate335(.out(and335), .in0(sizeov_not), .in1(modrm5), .in2(modrm4), .in3(modrm3), .in4(op15), .in5(op14), .in6(op13_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate336(.out(and336), .in0(modrm5
), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate337(.out(and337), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and5$ and_gate338(.out(and338), .in0(op15_not), .in1(op14), .in2(op13_not), .in3(op12), .in4(op11));
and5$ and_gate339(.out(and339), .in0(op15), .in1(op14_not), .in2(op13), .in3(op12), .in4(op11));
and5$ and_gate340(.out(and340), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and16$ and_gate341(.out(and341), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5
), .in12(op3), .in13(op2), .in14(op1), .in15(op0_not));
and16$ and_gate342(.out(and342), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7
), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate343(.out(and343), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op1), .in15(op0_not));
and17$ and_gate344(.out(and344), .in0(sizeov_not), .in1(op15
), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and11$ and_gate345(.out(and345), .in0(modrm5_not), .in1(modrm4), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13), .in6(op12), .in7(op11_not), .in8(op10
), .in9(op9), .in10(op8));
and16$ and_gate346(.out(and346), .in0(sizeov_not), .in1(op15_not), .in2(op14), .in3(op13), .in4(op12), .in5(op11_not), .in6(op10), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and15$ and_gate347(.out(and347), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13_not), .in4(op12_not), .in5(op10_not), .in6(op9), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate348(.out(and348), .in0(op15_not), .in1(op14_not), .in2(op13
), .in3(op12_not), .in4(op11_not), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and15$ and_gate349(.out(and349), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13), .in4(op12_not), .in5(op11_not), .in6(op9_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate350(.out(and350), .in0(op15_not), .in1(op14_not), .in2(op13), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate351(.out(and351), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate352(.out(and352), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2), .in15(op0));
and11$ and_gate353(.out(and353), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13), .in7(op12), .in8(op11_not), .in9(op10), .in10(op9));
and12$ and_gate354(.out(and354), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13), .in7(op12), .in8(op11
), .in9(op10), .in10(op9), .in11(op8));
and16$ and_gate355(.out(and355), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate356(.out(and356), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate357(.out(and357), .in0(sizeov_not), .in1(op15), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate358(.out(and358), .in0(modrm5), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op9_not), .in10(op8));
and11$ and_gate359(.out(and359), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and11$ and_gate360(.out(and360), .in0(sizeov_not), .in1(modrm5), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op8));
and5$ and_gate361(.out(and361), .in0(op15), .in1(op14_not), .in2(op13_not), .in3(op12), .in4(op11));
and17$ and_gate362(.out(and362), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5
), .in12(op4), .in13(op3), .in14(op2), .in15(op1_not), .in16(op0));
and16$ and_gate363(.out(and363), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8
), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3), .in13(op2), .in14(op1_not), .in15(op0_not));
and16$ and_gate364(.out(and364), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6), .in11(op5), .in12(op4_not), .in13(op3), .in14(op1), .in15(op0_not));
and17$ and_gate365(.out(and365), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13), .in4(op12_not), .in5(op11_not), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and11$ and_gate366(.out(and366), .in0(modrm5_not), .in1(modrm4), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13), .in6(op12), .in7(op11_not), .in8(op10), .in9(op9), .in10(op8));
and15$ and_gate367(.out(and367), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op9_not), .in6(op8), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and11$ and_gate368(.out(and368), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4), .in3(modrm3_not), .in4(op15), .in5(op14), .in6(op13), .in7(op12), .in8(op11_not), .in9(op10), .in10(op9));
and15$ and_gate369(.out(and369), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op9_not), .in7(op7_not), .in8(op6_not), .in9(op5_not), .in10(op4_not), .in11(op3_not), .in12(op2_not), .in13(op1_not), .in14(op0_not));
and16$ and_gate370(.out(and370), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11_not), .in5(op10_not), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate371(.out(and371), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11_not), .in6(op10_not), .in7(op9), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate372(.out(and372), .in0(sizeov_not), .in1(modrm5_not), .in2(modrm4_not), .in3(modrm3_not), .in4(op15), .in5(op14_not), .in6(op13_not), .in7(op12_not), .in8(op11_not), .in9(op10_not), .in10(op9_not));
and10$ and_gate373(.out(and373), .in0(modrm5), .in1(modrm4
), .in2(modrm3), .in3(op15), .in4(op14), .in5(op13_not), .in6(op12), .in7(op11_not), .in8(op10_not), .in9(op8));
and10$ and_gate374(.out(and374), .in0(sizeov_not), .in1(modrm5
), .in2(modrm4), .in3(modrm3), .in4(op15), .in5(op14), .in6(op13_not), .in7(op12), .in8(op11_not), .in9(op10_not));
and10$ and_gate375(.out(and375), .in0(modrm5), .in1(modrm4
), .in2(modrm3), .in3(op15), .in4(op14), .in5(op13_not), .in6(op11_not), .in7(op10_not), .in8(op9_not), .in9(op8));
and10$ and_gate376(.out(and376), .in0(sizeov_not), .in1(modrm5
), .in2(modrm4), .in3(modrm3), .in4(op15), .in5(op14), .in6(op13_not), .in7(op11_not), .in8(op10_not), .in9(op9_not));
and10$ and_gate377(.out(and377), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11_not), .in8(op10_not), .in9(op8));
and16$ and_gate378(.out(and378), .in0(op15_not), .in1(op14_not), .in2(op13_not), .in3(op12_not), .in4(op11), .in5(op10), .in6(op9), .in7(op8), .in8(op7), .in9(op6_not), .in10(op5), .in11(op4), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and16$ and_gate379(.out(and379), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8
), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4), .in13(op3_not), .in14(op2_not), .in15(op1_not));
and16$ and_gate380(.out(and380), .in0(sizeov_not), .in1(op15_not), .in2(op14), .in3(op13), .in4(op12
), .in5(op11_not), .in6(op10), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate381(.out(and381), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2), .in15(op0));
and16$ and_gate382(.out(and382), .in0(sizeov_not), .in1(op15_not), .in2(op14), .in3(op13), .in4(op12), .in5(op11_not), .in6(op10), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate383(.out(and383), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10
), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1), .in16(op0_not));
and16$ and_gate384(.out(and384), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2), .in15(op0));
and17$ and_gate385(.out(and385), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2), .in15(op1), .in16(op0));
and17$ and_gate386(.out(and386), .in0(sizeov_not), .in1(op15_not), .in2(op14), .in3(op13), .in4(op12), .in5(op11_not), .in6(op10
), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate387(.out(and387), .in0(sizeov_not), .in1(op15), .in2(op14), .in3(op13_not), .in4(op12_not), .in5(op10_not), .in6(op9), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate388(.out(and388), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11
), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op2_not), .in14(op1_not), .in15(op0));
and17$ and_gate389(.out(and389), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate390(.out(and390), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op11_not), .in5(op10), .in6(op9), .in7(op8), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate391(.out(and391), .in0(modrm5_not), .in1(modrm4_not), .in2(modrm3_not), .in3(op15), .in4(op14_not), .in5(op13_not), .in6(op12_not), .in7(op11), .in8(op10), .in9(op9), .in10(op8));
and5$ and_gate392(.out(and392), .in0(op15_not), .in1(op14), .in2(op13_not), .in3(op12), .in4(op11));
and16$ and_gate393(.out(and393), .in0(sizeov_not), .in1(op15_not), .in2(op14), .in3(op13), .in4(op12_not), .in5(op11), .in6(op10_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate394(.out(and394), .in0(op15_not), .in1(op14), .in2(op13), .in3(op12_not), .in4(op11), .in5(op10_not), .in6(op9_not), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and16$ and_gate395(.out(and395), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8), .in9(op7), .in10(op6_not), .in11(op5), .in12(op4_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and17$ and_gate396(.out(and396), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op12_not), .in5(op11), .in6(op10), .in7(op9), .in8(op8_not), .in9(op7_not), .in10(op6_not), .in11(op5_not), .in12(op4_not), .in13(op3_not), .in14(op2_not), .in15(op1_not), .in16(op0_not));
and16$ and_gate397(.out(and397), .in0(sizeov_not), .in1(op15_not), .in2(op14_not), .in3(op13_not), .in4(op11_not), .in5(op10), .in6(op9), .in7(op8_not), .in8(op7_not), .in9(op6_not), .in10(op5_not), .in11(op4_not), .in12(op3_not), .in13(op2_not), .in14(op1_not), .in15(op0_not));
and11$ and_gate398(.out(and398), .in0(modrm5), .in1(modrm4), .in2(modrm3_not), .in3(op15), .in4(op14), .in5(op13), .in6(op12), .in7(op11), .in8(op10), .in9(op9), .in10(op8));
and5$ and_gate399(.out(and399), .in0(op15_not), .in1(op14), .in2(op13_not), .in3(op12), .in4(op11));

or6$ or_gate0(.out(or0), .in0(and2), .in1(and3), .in2(and4), .in3(and5), .in4(and6), .in5(and7));
or43$ or_gate1(.out(or1), .in0(and8), .in1(and9), .in2(and10), .in3(and11), .in4(and12), .in5(and13), .in6(and14), .in7(and15), .in8(and16), .in9(and17), .in10(and18), .in11(and19), .in12(and20), .in13(and21), .in14(and22), .in15(and23), .in16(and24), .in17(and25), .in18(and26), .in19(and27), .in20(and28), .in21(and29), .in22(and30), .in23(and31), .in24(and32), .in25(and33), .in26(and34), .in27(and35), .in28(and36), .in29(and37), .in30(and38), .in31(and39), .in32(and40), .in33(and41), .in34(and42), .in35(and43), .in36(and44), .in37(and45), .in38(and46), .in39(and47), .in40(and48), .in41(and49), .in42(and50));
or37$ or_gate2(.out(or2), .in0(and51), .in1(and52), .in2(and53), .in3(and54), .in4(and55), .in5(and56), .in6(and57), .in7(and58), .in8(and59), .in9(and60), .in10(and61), .in11(and62), .in12(and63), .in13(and64), .in14(and65), .in15(and66), .in16(and67), .in17(and68), .in18(and69), .in19(and70), .in20(and71), .in21(and72), .in22(and73), .in23(and74), .in24(and75), .in25(and76), .in26(and77), .in27(and78), .in28(and79), .in29(and80), .in30(and81), .in31(and82), .in32(and83), .in33(and84), .in34(and85), .in35(and86), .in36(and87));
or37$ or_gate3(.out(or3), .in0(and88), .in1(and89), .in2(and90), .in3(and91), .in4(and92), .in5(and93), .in6(and94), .in7(and95), .in8(and96), .in9(and97), .in10(and98), .in11(and99), .in12(and100), .in13(and101), .in14(and102), .in15(and103), .in16(and104), .in17(and105), .in18(and106), .in19(and107), .in20(and108), .in21(and109), .in22(and110), .in23(and111), .in24(and112), .in25(and113), .in26(and114), .in27(and115), .in28(and116), .in29(and117), .in30(and118), .in31(and119), .in32(and120), .in33(and121), .in34(and122), .in35(and123), .in36(and124));
or9$ or_gate4(.out(or4), .in0(and125), .in1(and126), .in2(and127), .in3(and128), .in4(and129), .in5(and130), .in6(and131), .in7(and132), .in8(and133));
or26$ or_gate5(.out(or5), .in0(and134), .in1(and135), .in2(and136), .in3(and137), .in4(and138), .in5(and139), .in6(and140), .in7(and141), .in8(and142), .in9(and143), .in10(and144), .in11(and145), .in12(and146), .in13(and147), .in14(and148), .in15(and149), .in16(and150), .in17(and151), .in18(and152), .in19(and153), .in20(and154), .in21(and155), .in22(and156), .in23(and157), .in24(and158), .in25(and159));
or36$ or_gate6(.out(or6), .in0(and160), .in1(and161), .in2(and162), .in3(and163), .in4(and164), .in5(and165), .in6(and166), .in7(and167), .in8(and168), .in9(and169), .in10(and170), .in11(and171), .in12(and172), .in13(and173), .in14(and174), .in15(and175), .in16(and176), .in17(and177), .in18(and178), .in19(and179), .in20(and180), .in21(and181), .in22(and182), .in23(and183), .in24(and184), .in25(and185), .in26(and186), .in27(and187), .in28(and188), .in29(and189), .in30(and190), .in31(and191), .in32(and192), .in33(and193), .in34(and194), .in35(and195));
or6$ or_gate7(.out(or7), .in0(and196), .in1(and197), .in2(and198), .in3(and199), .in4(and200), .in5(and201));
or35$ or_gate8(.out(or8), .in0(and202), .in1(and203), .in2(and204), .in3(and205), .in4(and206), .in5(and207), .in6(and208), .in7(and209), .in8(and210), .in9(and211), .in10(and212), .in11(and213), .in12(and214), .in13(and215), .in14(and216), .in15(and217), .in16(and218), .in17(and219), .in18(and220), .in19(and221), .in20(and222), .in21(and223), .in22(and224), .in23(and225), .in24(and226), .in25(and227), .in26(and228), .in27(and229), .in28(and230), .in29(and231), .in30(and232), .in31(and233), .in32(and234), .in33(and235), .in34(and236));
or2$ or_gate9(.out(or9), .in0(and237), .in1(and238));
or15$ or_gate10(.out(or10), .in0(and239), .in1(and240), .in2(and241), .in3(and242), .in4(and243), .in5(and244), .in6(and245), .in7(and246), .in8(and247), .in9(and248), .in10(and249), .in11(and250), .in12(and251), .in13(and252), .in14(and253));
or2$ or_gate11(.out(or11), .in0(and254), .in1(and255));
or3$ or_gate12(.out(or12), .in0(and256), .in1(and257), .in2(and258));
or3$ or_gate13(.out(or13), .in0(and259), .in1(and260), .in2(and261));
or10$ or_gate14(.out(or14), .in0(and263), .in1(and264), .in2(and265), .in3(and266), .in4(and267), .in5(and268), .in6(and269), .in7(and270), .in8(and271), .in9(and272));
or4$ or_gate15(.out(or15), .in0(and273), .in1(and274), .in2(and275), .in3(and276));
or20$ or_gate16(.out(or16), .in0(and277), .in1(and278), .in2(and279), .in3(and280), .in4(and281), .in5(and282), .in6(and283), .in7(and284), .in8(and285), .in9(and286), .in10(and287), .in11(and288), .in12(and289), .in13(and290), .in14(and291), .in15(and292), .in16(and293), .in17(and294), .in18(and295), .in19(and296));
or44$ or_gate17(.out(or17), .in0(and297), .in1(and298), .in2(and299), .in3(and300), .in4(and301), .in5(and302), .in6(and303), .in7(and304), .in8(and305), .in9(and306), .in10(and307), .in11(and308), .in12(and309), .in13(and310), .in14(and311), .in15(and312), .in16(and313), .in17(and314), .in18(and315), .in19(and316), .in20(and317), .in21(and318), .in22(and319), .in23(and320), .in24(and321), .in25(and322), .in26(and323), .in27(and324), .in28(and325), .in29(and326), .in30(and327), .in31(and328), .in32(and329), .in33(and330), .in34(and331), .in35(and332), .in36(and333), .in37(and334), .in38(and335), .in39(and336), .in40(and337), .in41(and338), .in42(and339), .in43(and340));
or21$ or_gate18(.out(or18), .in0(and341), .in1(and342), .in2(and343), .in3(and344), .in4(and345), .in5(and346), .in6(and347), .in7(and348), .in8(and349), .in9(and350), .in10(and351), .in11(and352), .in12(and353), .in13(and354), .in14(and355), .in15(and356), .in16(and357), .in17(and358), .in18(and359), .in19(and360), .in20(and361));
or16$ or_gate19(.out(or19), .in0(and362), .in1(and363), .in2(and364), .in3(and365), .in4(and366), .in5(and367), .in6(and368), .in7(and369), .in8(and370), .in9(and371), .in10(and372), .in11(and373), .in12(and374), .in13(and375), .in14(and376), .in15(and377));
or4$ or_gate20(.out(or20), .in0(and378), .in1(and379), .in2(and380), .in3(and381));
or3$ or_gate21(.out(or21), .in0(and382), .in1(and383), .in2(and384));
or2$ or_gate22(.out(or22), .in0(and385), .in1(and386));
or6$ or_gate23(.out(or23), .in0(and387), .in1(and388), .in2(and389), .in3(and390), .in4(and391), .in5(and392));
or7$ or_gate24(.out(or24), .in0(and393), .in1(and394), .in2(and395), .in3(and396), .in4(and397), .in5(and398), .in6(and399));

assign setd = and0;
assign cleard = and1;
assign size2 = or0;
assign size1 = or1;
assign size0 = or2;
assign op0_2 = or3;
assign op0_1 = or4;
assign op0_0 = or5;
assign op1_2 = or6;
assign op1_1 = or7;
assign op1_0 = or8;
assign op0_reg_4 = or9;
assign op0_reg_3 = or10;
assign op0_reg_2 = or11;
assign op0_reg_1 = or12;
assign op0_reg_0 = or13;
assign op1_reg_4 = and262;
assign op1_reg_3 = or14;
assign op1_reg_2 = or14;
assign op1_reg_1 = or14;
assign op1_reg_0 = or15;
assign alu_op_3 = or16;
assign alu_op_2 = or17;
assign alu_op_1 = or18;
assign alu_op_0 = or19;
assign flag0_2 = or19;
assign flag0_1 = or20;
assign flag0_0 = or21;
assign flag1_2 = or21;
assign flag1_1 = or21;
assign flag1_0 = or22;
assign stack_op_1 = or23;
assign stack_op_0 = or24;

endmodule
