`timescale 1ns/1ps
/*//and$ modules larger than 4 inputs
module and5$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4);


wire AND0, AND1, AND_OUT;

and3$ g_and0(.in0(in0), .in1(in1), .in2(in2), .out(AND0));
and2$ g_and1(.in0(in3), .in1(in4), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and6$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5);


wire AND0, AND1, AND_OUT;

and3$ g_and0(.in0(in0), .in1(in1), .in2(in2), .out(AND0));
and3$ g_and1(.in0(in3), .in1(in4), .in2(in5), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and7$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6);


wire AND0, AND1, AND_OUT;

and3$ g_and0(.in0(in0), .in1(in1), .in2(in2), .out(AND0));
and4$ g_and1(.in0(in3), .in1(in4), .in2(in5), .in3(in6), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and8$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7);


wire AND0, AND1, AND_OUT;

and4$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .out(AND0));
and4$ g_and1(.in0(in4), .in1(in5), .in2(in6), .in3(in7), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and9$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8);


wire AND0, AND1, AND_OUT;

and4$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .out(AND0));
and5$ g_and1(.in0(in4), .in1(in5), .in2(in6), .in3(in7), .in4(in8), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and10$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9);


wire AND0, AND1, AND_OUT;

and5$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .out(AND0));
and5$ g_and1(.in0(in5), .in1(in6), .in2(in7), .in3(in8), .in4(in9), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and11$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10);


wire AND0, AND1, AND_OUT;

and5$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .out(AND0));
and6$ g_and1(.in0(in5), .in1(in6), .in2(in7), .in3(in8), .in4(in9), .in5(in10), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and12$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11);


wire AND0, AND1, AND_OUT;

and6$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .out(AND0));
and6$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and13$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12);


wire AND0, AND1, AND_OUT;

and6$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .out(AND0));
and7$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and14$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13);


wire AND0, AND1, AND_OUT;

and7$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .out(AND0));
and7$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and15$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14);


wire AND0, AND1, AND_OUT;

and7$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .out(AND0));
and8$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and16$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15);


wire AND0, AND1, AND_OUT;

and8$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .out(AND0));
and8$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and17$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16);


wire AND0, AND1, AND_OUT;

and8$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .out(AND0));
and9$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and18$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17);


wire AND0, AND1, AND_OUT;

and9$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .out(AND0));
and9$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and19$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18);


wire AND0, AND1, AND_OUT;

and9$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .out(AND0));
and10$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and20$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18,
input in19);


wire AND0, AND1, AND_OUT;

and10$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .in9(in19), .out(AND0));
and10$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and21$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18,
input in19,
input in20);


wire AND0, AND1, AND_OUT;

and10$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .in9(in19), .out(AND0));
and11$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .in10(in20), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));
endmodule

`timescale 1ns / 1ps
module and22$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18,
input in19,
input in20,
input in21);


wire AND0, AND1, AND_OUT;

and11$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .in9(in19), .in10(in21), .out(AND0));
and11$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .in10(in20), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and23$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18,
input in19,
input in20,
input in21,
input in22);


wire AND0, AND1, AND_OUT;

and11$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .in9(in19), .in10(in21), .out(AND0));
and12$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .in10(in20), .in11(in22), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and24$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18,
input in19,
input in20,
input in21,
input in22,
input in23);


wire AND0, AND1, AND_OUT;

and12$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .in9(in19), .in10(in21), .in11(in23), .out(AND0));
and12$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .in10(in20), .in11(in22), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule
*/
`timescale 1ns / 1ps
module and25$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18,
input in19,
input in20,
input in21,
input in22,
input in23,
input in24);


wire AND0, AND1, AND_OUT;

and12$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .in9(in19), .in10(in21), .in11(in23), .out(AND0));
and13$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .in10(in20), .in11(in22), .in12(in24), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and26$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18,
input in19,
input in20,
input in21,
input in22,
input in23,
input in24,
input in25);


wire AND0, AND1, AND_OUT;

and13$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .in9(in19), .in10(in21), .in11(in23), .in12(in25), .out(AND0));
and13$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .in10(in20), .in11(in22), .in12(in24), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and27$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18,
input in19,
input in20,
input in21,
input in22,
input in23,
input in24,
input in25,
input in26);


wire AND0, AND1, AND_OUT;

and13$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .in9(in19), .in10(in21), .in11(in23), .in12(in25), .out(AND0));
and14$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .in10(in20), .in11(in22), .in12(in24), .in13(in26), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and28$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18,
input in19,
input in20,
input in21,
input in22,
input in23,
input in24,
input in25,
input in26,
input in27);


wire AND0, AND1, AND_OUT;

and14$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .in9(in19), .in10(in21), .in11(in23), .in12(in25), .in13(in27), .out(AND0));
and14$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .in10(in20), .in11(in22), .in12(in24), .in13(in26), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and29$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18,
input in19,
input in20,
input in21,
input in22,
input in23,
input in24,
input in25,
input in26,
input in27,
input in28);


wire AND0, AND1, AND_OUT;

and14$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .in9(in19), .in10(in21), .in11(in23), .in12(in25), .in13(in27), .out(AND0));
and15$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .in10(in20), .in11(in22), .in12(in24), .in13(in26), .in14(in28), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and30$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18,
input in19,
input in20,
input in21,
input in22,
input in23,
input in24,
input in25,
input in26,
input in27,
input in28,
input in29);


wire AND0, AND1, AND_OUT;

and15$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .in9(in19), .in10(in21), .in11(in23), .in12(in25), .in13(in27), .in14(in29), .out(AND0));
and15$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .in10(in20), .in11(in22), .in12(in24), .in13(in26), .in14(in28), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and31$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18,
input in19,
input in20,
input in21,
input in22,
input in23,
input in24,
input in25,
input in26,
input in27,
input in28,
input in29,
input in30);


wire AND0, AND1, AND_OUT;

and15$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .in9(in19), .in10(in21), .in11(in23), .in12(in25), .in13(in27), .in14(in29), .out(AND0));
and16$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .in10(in20), .in11(in22), .in12(in24), .in13(in26), .in14(in28), .in15(in30), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule

`timescale 1ns / 1ps
module and32$(output out,
input in0, 
input in1, 
input in2, 
input in3, 
input in4,
input in5,
input in6,
input in7,
input in8,
input in9,
input in10,
input in11,
input in12,
input in13,
input in14,
input in15,
input in16,
input in17,
input in18,
input in19,
input in20,
input in21,
input in22,
input in23,
input in24,
input in25,
input in26,
input in27,
input in28,
input in29,
input in30,
input in31);


wire AND0, AND1, AND_OUT;

and16$ g_and0(.in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in13), .in7(in15), .in8(in17), .in9(in19), .in10(in21), .in11(in23), .in12(in25), .in13(in27), .in14(in29), .in15(in31), .out(AND0));
and16$ g_and1(.in0(in6), .in1(in7), .in2(in8), .in3(in9), .in4(in10), .in5(in11), .in6(in12), .in7(in14), .in8(in16), .in9(in18), .in10(in20), .in11(in22), .in12(in24), .in13(in26), .in14(in28), .in15(in30), .out(AND1));
and2$ g_and_out(.in0(AND0), .in1(AND1), .out(out));

endmodule